* Extracted by KLayout with SG13G2 LVS runset on : 29/04/2024 05:18

* cell sg13g2_Clamp_N20N0D
* pin pad
* pin iovss
.SUBCKT sg13g2_Clamp_N20N0D pad iovss
* device instance $1 r0 *1 25.52,4.95 sg13_hv_nmos
M$1 iovss \$5 pad iovss sg13_hv_nmos W=88.00000000000001 L=0.5999999999999998
* device instance $21 r0 *1 66.305,2.75 res_rppd
R$21 iovss \$5 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0 ps=0.0
+ m=1.0
.ENDS sg13g2_Clamp_N20N0D

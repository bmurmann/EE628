* Extracted by KLayout with SG13G2 LVS runset on : 03/05/2024 05:38

* cell sg13g2_Clamp_N43N43D4R
* pin sub!
.SUBCKT sg13g2_Clamp_N43N43D4R sub!
* device instance $1 r0 *1 8.155,4.95 sg13_hv_nmos
M$1 sub! \$5 \$6 sub! sg13_hv_nmos W=756.7999999999977 L=0.5999999999999998
* device instance $173 r0 *1 4.765,21.35 dantenna
D$173 sub! \$5 dantenna A=0.192 P=1.88 m=1
.ENDS sg13g2_Clamp_N43N43D4R

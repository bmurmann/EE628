* Extracted by KLayout with SG13G2 LVS runset on : 03/05/2024 20:54

* cell padring
* pin PAD,RES
* pin CK4,PAD
* pin CK5,PAD
* pin CK6,PAD
* pin IOVDD
* pin AVDD
* pin CORE
* pin CORE
* pin VDD
* pin CORE
* pin CORE
* pin res_c
* pin ck4_c
* pin ck5_c
* pin ck6_c
* pin IN6,PAD
* pin OUT6
* pin out6_c
* pin CORE,in6_c
* pin IN5,PAD
* pin OUT5
* pin out5_c
* pin CORE,in5_c
* pin IN4,PAD
* pin OUT4
* pin out4_c
* pin CORE,in4_c
* pin PAD,VLO
* pin CORE
* pin PAD,VHI
* pin CORE
* pin IN3,PAD
* pin OUT3
* pin out3_c
* pin CORE,in3_c
* pin IN2,PAD
* pin OUT2
* pin out2_c
* pin CORE,in2_c
* pin IN1,PAD
* pin OUT1
* pin out1_c
* pin CORE,in1_c
* pin PAD,VREF
* pin CORE,vref_c
* pin PAD,VLDO
* pin ck3_c
* pin ck2_c
* pin ck1_c
* pin CORE
* pin CORE
* pin CORE
* pin CORE
* pin CK3,PAD
* pin CK2,PAD
* pin CK1,PAD
* pin VSS
.SUBCKT padring PAD|RES CK4|PAD CK5|PAD CK6|PAD IOVDD AVDD CORE CORE$1 VDD
+ CORE$2 CORE$3 res_c ck4_c ck5_c ck6_c IN6|PAD OUT6 out6_c CORE|in6_c IN5|PAD
+ OUT5 out5_c CORE|in5_c IN4|PAD OUT4 out4_c CORE|in4_c PAD|VLO CORE$4 PAD|VHI
+ CORE$5 IN3|PAD OUT3 out3_c CORE|in3_c IN2|PAD OUT2 out2_c CORE|in2_c IN1|PAD
+ OUT1 out1_c CORE|in1_c PAD|VREF CORE|vref_c PAD|VLDO ck3_c ck2_c ck1_c CORE$6
+ CORE$7 CORE$8 CORE$9 CK3|PAD CK2|PAD CK1|PAD VSS
* device instance $1 r0 *1 240.255,159.005 sg13_lv_nmos
M$1 res_c \$178 VSS VSS sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $2 r0 *1 440.255,159.005 sg13_lv_nmos
M$2 ck4_c \$179 VSS VSS sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $3 r0 *1 540.255,159.005 sg13_lv_nmos
M$3 ck5_c \$180 VSS VSS sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $4 r0 *1 640.255,159.005 sg13_lv_nmos
M$4 ck6_c \$181 VSS VSS sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $5 r0 *1 800.995,217.48 sg13_lv_nmos
M$5 \$227 out6_c VSS VSS sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $6 r0 *1 800.995,220.99 sg13_lv_nmos
M$6 \$255 out6_c VSS VSS sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $7 r0 *1 800.995,317.48 sg13_lv_nmos
M$7 \$340 out5_c VSS VSS sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $8 r0 *1 800.995,320.99 sg13_lv_nmos
M$8 \$368 out5_c VSS VSS sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $9 r0 *1 800.995,417.48 sg13_lv_nmos
M$9 \$453 out4_c VSS VSS sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $10 r0 *1 800.995,420.99 sg13_lv_nmos
M$10 \$481 out4_c VSS VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $11 r0 *1 800.995,717.48 sg13_lv_nmos
M$11 \$714 out3_c VSS VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $12 r0 *1 800.995,720.99 sg13_lv_nmos
M$12 \$742 out3_c VSS VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $13 r0 *1 800.995,817.48 sg13_lv_nmos
M$13 \$827 out2_c VSS VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $14 r0 *1 800.995,820.99 sg13_lv_nmos
M$14 \$855 out2_c VSS VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $15 r0 *1 800.995,917.48 sg13_lv_nmos
M$15 \$940 out1_c VSS VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $16 r0 *1 800.995,920.99 sg13_lv_nmos
M$16 \$968 out1_c VSS VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $17 r0 *1 440.255,980.995 sg13_lv_nmos
M$17 ck3_c \$1036 VSS VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $18 r0 *1 540.255,980.995 sg13_lv_nmos
M$18 ck2_c \$1037 VSS VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $19 r0 *1 640.255,980.995 sg13_lv_nmos
M$19 ck1_c \$1038 VSS VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $20 r0 *1 241.765,159.055 sg13_hv_nmos
M$20 VSS CORE \$178 VSS sg13_hv_nmos W=2.6499999999999995 L=0.4499999999999999
* device instance $21 r0 *1 441.765,159.055 sg13_hv_nmos
M$21 VSS CORE$1 \$179 VSS sg13_hv_nmos W=2.6499999999999995 L=0.4499999999999999
* device instance $22 r0 *1 541.765,159.055 sg13_hv_nmos
M$22 VSS CORE$2 \$180 VSS sg13_hv_nmos W=2.6499999999999995 L=0.4499999999999999
* device instance $23 r0 *1 641.765,159.055 sg13_hv_nmos
M$23 VSS CORE$3 \$181 VSS sg13_hv_nmos W=2.6499999999999995 L=0.4499999999999999
* device instance $24 r0 *1 -169.05,205.52 sg13_hv_nmos
M$24 VSS \$217 IN6|PAD VSS sg13_hv_nmos W=88.00000000000001 L=0.5999999999999998
* device instance $44 r0 *1 949.05,214.58 sg13_hv_nmos
M$44 VSS \$244 OUT6 VSS sg13_hv_nmos W=35.199999999999996 L=0.5999999999999998
* device instance $52 r0 *1 804.68,217.64 sg13_hv_nmos
M$52 \$228 out6_c VSS VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $53 r0 *1 804.68,218.47 sg13_hv_nmos
M$53 VSS \$227 \$238 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $54 r0 *1 804.68,219.81 sg13_hv_nmos
M$54 VSS \$238 \$244 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $55 r0 *1 804.68,221.15 sg13_hv_nmos
M$55 \$256 out6_c VSS VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $56 r0 *1 804.68,221.98 sg13_hv_nmos
M$56 VSS \$255 \$263 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $57 r0 *1 804.68,223.32 sg13_hv_nmos
M$57 VSS \$263 \$208 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $58 r0 *1 -169.05,305.52 sg13_hv_nmos
M$58 VSS \$330 IN5|PAD VSS sg13_hv_nmos W=88.00000000000001 L=0.5999999999999998
* device instance $78 r0 *1 949.05,314.58 sg13_hv_nmos
M$78 VSS \$357 OUT5 VSS sg13_hv_nmos W=35.199999999999996 L=0.5999999999999998
* device instance $86 r0 *1 804.68,317.64 sg13_hv_nmos
M$86 \$341 out5_c VSS VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $87 r0 *1 804.68,318.47 sg13_hv_nmos
M$87 VSS \$340 \$351 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $88 r0 *1 804.68,319.81 sg13_hv_nmos
M$88 VSS \$351 \$357 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $89 r0 *1 804.68,321.15 sg13_hv_nmos
M$89 \$369 out5_c VSS VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $90 r0 *1 804.68,321.98 sg13_hv_nmos
M$90 VSS \$368 \$376 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $91 r0 *1 804.68,323.32 sg13_hv_nmos
M$91 VSS \$376 \$321 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $92 r0 *1 -169.05,405.52 sg13_hv_nmos
M$92 VSS \$443 IN4|PAD VSS sg13_hv_nmos W=88.00000000000001 L=0.5999999999999998
* device instance $112 r0 *1 949.05,414.58 sg13_hv_nmos
M$112 VSS \$470 OUT4 VSS sg13_hv_nmos W=35.199999999999996 L=0.5999999999999998
* device instance $120 r0 *1 804.68,417.64 sg13_hv_nmos
M$120 \$454 out4_c VSS VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $121 r0 *1 804.68,418.47 sg13_hv_nmos
M$121 VSS \$453 \$464 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $122 r0 *1 804.68,419.81 sg13_hv_nmos
M$122 VSS \$464 \$470 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $123 r0 *1 804.68,421.15 sg13_hv_nmos
M$123 \$482 out4_c VSS VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $124 r0 *1 804.68,421.98 sg13_hv_nmos
M$124 VSS \$481 \$489 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $125 r0 *1 804.68,423.32 sg13_hv_nmos
M$125 VSS \$489 \$434 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $126 r0 *1 -169.05,505.52 sg13_hv_nmos
M$126 VSS \$559 PAD|VLO VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $146 r0 *1 879.21,583.22 sg13_hv_nmos
M$146 VSS \$620 \$619 VSS sg13_hv_nmos W=107.99999999999999 L=0.4999999999999999
* device instance $152 r0 *1 879.21,593 sg13_hv_nmos
M$152 VSS \$620 VSS VSS sg13_hv_nmos W=125.99999999999999 L=9.499999999999996
* device instance $172 r0 *1 934.53,588.155 sg13_hv_nmos
M$172 VSS \$619 IOVDD VSS sg13_hv_nmos W=756.7999999999977 L=0.5999999999999998
* device instance $344 r0 *1 -169.05,605.52 sg13_hv_nmos
M$344 VSS \$625 PAD|VHI VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $364 r0 *1 -169.05,705.52 sg13_hv_nmos
M$364 VSS \$704 IN3|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $384 r0 *1 949.05,714.58 sg13_hv_nmos
M$384 VSS \$731 OUT3 VSS sg13_hv_nmos W=35.199999999999996 L=0.5999999999999998
* device instance $392 r0 *1 804.68,717.64 sg13_hv_nmos
M$392 \$715 out3_c VSS VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $393 r0 *1 804.68,718.47 sg13_hv_nmos
M$393 VSS \$714 \$725 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $394 r0 *1 804.68,719.81 sg13_hv_nmos
M$394 VSS \$725 \$731 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $395 r0 *1 804.68,721.15 sg13_hv_nmos
M$395 \$743 out3_c VSS VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $396 r0 *1 804.68,721.98 sg13_hv_nmos
M$396 VSS \$742 \$750 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $397 r0 *1 804.68,723.32 sg13_hv_nmos
M$397 VSS \$750 \$695 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $398 r0 *1 -169.05,805.52 sg13_hv_nmos
M$398 VSS \$817 IN2|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $418 r0 *1 949.05,814.58 sg13_hv_nmos
M$418 VSS \$844 OUT2 VSS sg13_hv_nmos W=35.199999999999996 L=0.5999999999999998
* device instance $426 r0 *1 804.68,817.64 sg13_hv_nmos
M$426 \$828 out2_c VSS VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $427 r0 *1 804.68,818.47 sg13_hv_nmos
M$427 VSS \$827 \$838 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $428 r0 *1 804.68,819.81 sg13_hv_nmos
M$428 VSS \$838 \$844 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $429 r0 *1 804.68,821.15 sg13_hv_nmos
M$429 \$856 out2_c VSS VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $430 r0 *1 804.68,821.98 sg13_hv_nmos
M$430 VSS \$855 \$863 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $431 r0 *1 804.68,823.32 sg13_hv_nmos
M$431 VSS \$863 \$808 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $432 r0 *1 -169.05,905.52 sg13_hv_nmos
M$432 VSS \$930 IN1|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $452 r0 *1 949.05,914.58 sg13_hv_nmos
M$452 VSS \$957 OUT1 VSS sg13_hv_nmos W=35.199999999999996 L=0.5999999999999998
* device instance $460 r0 *1 804.68,917.64 sg13_hv_nmos
M$460 \$941 out1_c VSS VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $461 r0 *1 804.68,918.47 sg13_hv_nmos
M$461 VSS \$940 \$951 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $462 r0 *1 804.68,919.81 sg13_hv_nmos
M$462 VSS \$951 \$957 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $463 r0 *1 804.68,921.15 sg13_hv_nmos
M$463 \$969 out1_c VSS VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $464 r0 *1 804.68,921.98 sg13_hv_nmos
M$464 VSS \$968 \$976 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $465 r0 *1 804.68,923.32 sg13_hv_nmos
M$465 VSS \$976 \$921 VSS sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $466 r0 *1 441.765,980.945 sg13_hv_nmos
M$466 VSS CORE$6 \$1036 VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $467 r0 *1 541.765,980.945 sg13_hv_nmos
M$467 VSS CORE$7 \$1037 VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $468 r0 *1 641.765,980.945 sg13_hv_nmos
M$468 VSS CORE$8 \$1038 VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $469 r0 *1 3.22,1059.21 sg13_hv_nmos
M$469 VSS \$1164 \$1105 VSS sg13_hv_nmos W=107.99999999999999
+ L=0.4999999999999999
* device instance $475 r0 *1 13,1059.21 sg13_hv_nmos
M$475 VSS \$1164 VSS VSS sg13_hv_nmos W=125.99999999999999 L=9.499999999999996
* device instance $482 r0 *1 303.22,1059.21 sg13_hv_nmos
M$482 VSS \$1165 \$1106 VSS sg13_hv_nmos W=107.99999999999999
+ L=0.4999999999999999
* device instance $488 r0 *1 313,1059.21 sg13_hv_nmos
M$488 VSS \$1165 VSS VSS sg13_hv_nmos W=125.99999999999999 L=9.499999999999996
* device instance $495 r0 *1 703.22,1059.21 sg13_hv_nmos
M$495 VSS \$1166 \$1107 VSS sg13_hv_nmos W=107.99999999999999
+ L=0.4999999999999999
* device instance $501 r0 *1 713,1059.21 sg13_hv_nmos
M$501 VSS \$1166 VSS VSS sg13_hv_nmos W=125.99999999999999 L=9.499999999999996
* device instance $547 r0 *1 8.155,1114.53 sg13_hv_nmos
M$547 VSS \$1105 AVDD VSS sg13_hv_nmos W=756.7999999999977 L=0.5999999999999998
* device instance $590 r0 *1 308.155,1114.53 sg13_hv_nmos
M$590 VSS \$1106 IOVDD VSS sg13_hv_nmos W=756.7999999999977 L=0.5999999999999998
* device instance $633 r0 *1 708.155,1114.53 sg13_hv_nmos
M$633 VSS \$1107 VDD VSS sg13_hv_nmos W=756.7999999999977 L=0.5999999999999998
* device instance $977 r0 *1 125.52,1129.05 sg13_hv_nmos
M$977 VSS \$1236 PAD|VREF VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $997 r0 *1 225.52,1129.05 sg13_hv_nmos
M$997 VSS \$1237 PAD|VLDO VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $1103 r0 *1 240.255,163.995 sg13_lv_pmos
M$1103 res_c \$178 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1104 r0 *1 440.255,163.995 sg13_lv_pmos
M$1104 ck4_c \$179 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1105 r0 *1 540.255,163.995 sg13_lv_pmos
M$1105 ck5_c \$180 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1106 r0 *1 640.255,163.995 sg13_lv_pmos
M$1106 ck6_c \$181 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1107 r0 *1 796.005,217.48 sg13_lv_pmos
M$1107 \$227 out6_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1108 r0 *1 796.005,220.99 sg13_lv_pmos
M$1108 \$255 out6_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1109 r0 *1 796.005,317.48 sg13_lv_pmos
M$1109 \$340 out5_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1110 r0 *1 796.005,320.99 sg13_lv_pmos
M$1110 \$368 out5_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1111 r0 *1 796.005,417.48 sg13_lv_pmos
M$1111 \$453 out4_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1112 r0 *1 796.005,420.99 sg13_lv_pmos
M$1112 \$481 out4_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1113 r0 *1 796.005,717.48 sg13_lv_pmos
M$1113 \$714 out3_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1114 r0 *1 796.005,720.99 sg13_lv_pmos
M$1114 \$742 out3_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1115 r0 *1 796.005,817.48 sg13_lv_pmos
M$1115 \$827 out2_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1116 r0 *1 796.005,820.99 sg13_lv_pmos
M$1116 \$855 out2_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1117 r0 *1 796.005,917.48 sg13_lv_pmos
M$1117 \$940 out1_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1118 r0 *1 796.005,920.99 sg13_lv_pmos
M$1118 \$968 out1_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1119 r0 *1 440.255,976.005 sg13_lv_pmos
M$1119 ck3_c \$1036 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1120 r0 *1 540.255,976.005 sg13_lv_pmos
M$1120 ck2_c \$1037 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1121 r0 *1 640.255,976.005 sg13_lv_pmos
M$1121 ck1_c \$1038 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1122 r0 *1 241.765,163.945 sg13_hv_pmos
M$1122 VDD CORE \$178 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1123 r0 *1 441.765,163.945 sg13_hv_pmos
M$1123 VDD CORE$1 \$179 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1124 r0 *1 541.765,163.945 sg13_hv_pmos
M$1124 VDD CORE$2 \$180 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1125 r0 *1 641.765,163.945 sg13_hv_pmos
M$1125 VDD CORE$3 \$181 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1126 r0 *1 -108.92,205.52 sg13_hv_pmos
M$1126 AVDD \$218 IN6|PAD AVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1166 r0 *1 881.82,214.58 sg13_hv_pmos
M$1166 IOVDD \$208 OUT6 IOVDD sg13_hv_pmos W=106.55999999999996
+ L=0.5999999999999999
* device instance $1182 r0 *1 808.82,217.64 sg13_hv_pmos
M$1182 \$228 \$238 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1183 r0 *1 808.82,218.47 sg13_hv_pmos
M$1183 IOVDD \$228 \$238 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1184 r0 *1 808.82,219.81 sg13_hv_pmos
M$1184 IOVDD \$238 \$244 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1185 r0 *1 808.82,221.15 sg13_hv_pmos
M$1185 \$256 \$263 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1186 r0 *1 808.82,221.98 sg13_hv_pmos
M$1186 IOVDD \$256 \$263 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1187 r0 *1 808.82,223.32 sg13_hv_pmos
M$1187 IOVDD \$263 \$208 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1188 r0 *1 -108.92,305.52 sg13_hv_pmos
M$1188 AVDD \$331 IN5|PAD AVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1228 r0 *1 881.82,314.58 sg13_hv_pmos
M$1228 IOVDD \$321 OUT5 IOVDD sg13_hv_pmos W=106.55999999999996
+ L=0.5999999999999999
* device instance $1244 r0 *1 808.82,317.64 sg13_hv_pmos
M$1244 \$341 \$351 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1245 r0 *1 808.82,318.47 sg13_hv_pmos
M$1245 IOVDD \$341 \$351 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1246 r0 *1 808.82,319.81 sg13_hv_pmos
M$1246 IOVDD \$351 \$357 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1247 r0 *1 808.82,321.15 sg13_hv_pmos
M$1247 \$369 \$376 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1248 r0 *1 808.82,321.98 sg13_hv_pmos
M$1248 IOVDD \$369 \$376 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1249 r0 *1 808.82,323.32 sg13_hv_pmos
M$1249 IOVDD \$376 \$321 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1250 r0 *1 -108.92,405.52 sg13_hv_pmos
M$1250 AVDD \$444 IN4|PAD AVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1290 r0 *1 881.82,414.58 sg13_hv_pmos
M$1290 IOVDD \$434 OUT4 IOVDD sg13_hv_pmos W=106.55999999999996
+ L=0.5999999999999999
* device instance $1306 r0 *1 808.82,417.64 sg13_hv_pmos
M$1306 \$454 \$464 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1307 r0 *1 808.82,418.47 sg13_hv_pmos
M$1307 IOVDD \$454 \$464 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1308 r0 *1 808.82,419.81 sg13_hv_pmos
M$1308 IOVDD \$464 \$470 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1309 r0 *1 808.82,421.15 sg13_hv_pmos
M$1309 \$482 \$489 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1310 r0 *1 808.82,421.98 sg13_hv_pmos
M$1310 IOVDD \$482 \$489 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1311 r0 *1 808.82,423.32 sg13_hv_pmos
M$1311 IOVDD \$489 \$434 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1312 r0 *1 -108.92,505.52 sg13_hv_pmos
M$1312 AVDD \$560 PAD|VLO AVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1352 r0 *1 865.09,598.44 sg13_hv_pmos
M$1352 IOVDD \$620 \$619 IOVDD sg13_hv_pmos W=349.99999999999994
+ L=0.4999999999999999
* device instance $1402 r0 *1 -108.92,605.52 sg13_hv_pmos
M$1402 AVDD \$626 PAD|VHI AVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1442 r0 *1 -108.92,705.52 sg13_hv_pmos
M$1442 AVDD \$705 IN3|PAD AVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1482 r0 *1 881.82,714.58 sg13_hv_pmos
M$1482 IOVDD \$695 OUT3 IOVDD sg13_hv_pmos W=106.55999999999996
+ L=0.5999999999999999
* device instance $1498 r0 *1 808.82,717.64 sg13_hv_pmos
M$1498 \$715 \$725 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1499 r0 *1 808.82,718.47 sg13_hv_pmos
M$1499 IOVDD \$715 \$725 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1500 r0 *1 808.82,719.81 sg13_hv_pmos
M$1500 IOVDD \$725 \$731 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1501 r0 *1 808.82,721.15 sg13_hv_pmos
M$1501 \$743 \$750 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1502 r0 *1 808.82,721.98 sg13_hv_pmos
M$1502 IOVDD \$743 \$750 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1503 r0 *1 808.82,723.32 sg13_hv_pmos
M$1503 IOVDD \$750 \$695 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1504 r0 *1 -108.92,805.52 sg13_hv_pmos
M$1504 AVDD \$818 IN2|PAD AVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1544 r0 *1 881.82,814.58 sg13_hv_pmos
M$1544 IOVDD \$808 OUT2 IOVDD sg13_hv_pmos W=106.55999999999996
+ L=0.5999999999999999
* device instance $1560 r0 *1 808.82,817.64 sg13_hv_pmos
M$1560 \$828 \$838 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1561 r0 *1 808.82,818.47 sg13_hv_pmos
M$1561 IOVDD \$828 \$838 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1562 r0 *1 808.82,819.81 sg13_hv_pmos
M$1562 IOVDD \$838 \$844 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1563 r0 *1 808.82,821.15 sg13_hv_pmos
M$1563 \$856 \$863 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1564 r0 *1 808.82,821.98 sg13_hv_pmos
M$1564 IOVDD \$856 \$863 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1565 r0 *1 808.82,823.32 sg13_hv_pmos
M$1565 IOVDD \$863 \$808 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1566 r0 *1 -108.92,905.52 sg13_hv_pmos
M$1566 AVDD \$931 IN1|PAD AVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1606 r0 *1 881.82,914.58 sg13_hv_pmos
M$1606 IOVDD \$921 OUT1 IOVDD sg13_hv_pmos W=106.55999999999996
+ L=0.5999999999999999
* device instance $1622 r0 *1 808.82,917.64 sg13_hv_pmos
M$1622 \$941 \$951 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1623 r0 *1 808.82,918.47 sg13_hv_pmos
M$1623 IOVDD \$941 \$951 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1624 r0 *1 808.82,919.81 sg13_hv_pmos
M$1624 IOVDD \$951 \$957 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1625 r0 *1 808.82,921.15 sg13_hv_pmos
M$1625 \$969 \$976 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1626 r0 *1 808.82,921.98 sg13_hv_pmos
M$1626 IOVDD \$969 \$976 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1627 r0 *1 808.82,923.32 sg13_hv_pmos
M$1627 IOVDD \$976 \$921 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1628 r0 *1 441.765,976.055 sg13_hv_pmos
M$1628 VDD CORE$6 \$1036 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1629 r0 *1 541.765,976.055 sg13_hv_pmos
M$1629 VDD CORE$7 \$1037 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1630 r0 *1 641.765,976.055 sg13_hv_pmos
M$1630 VDD CORE$8 \$1038 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1631 r0 *1 18.44,1045.09 sg13_hv_pmos
M$1631 AVDD \$1164 \$1105 AVDD sg13_hv_pmos W=349.99999999999994
+ L=0.4999999999999999
* device instance $1681 r0 *1 318.44,1045.09 sg13_hv_pmos
M$1681 IOVDD \$1165 \$1106 IOVDD sg13_hv_pmos W=349.99999999999994
+ L=0.4999999999999999
* device instance $1731 r0 *1 718.44,1045.09 sg13_hv_pmos
M$1731 IOVDD \$1166 \$1107 IOVDD sg13_hv_pmos W=349.99999999999994
+ L=0.4999999999999999
* device instance $1781 r0 *1 125.52,1061.82 sg13_hv_pmos
M$1781 AVDD \$1122 PAD|VREF AVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1821 r0 *1 225.52,1061.82 sg13_hv_pmos
M$1821 AVDD \$1123 PAD|VLDO AVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1861 r0 *1 4.54,24.19 dantenna
D$1861 VSS VSS dantenna A=35.0028 P=58.08 m=10
* device instance $1865 r0 *1 204.54,24.19 dantenna
D$1865 VSS PAD|RES dantenna A=35.0028 P=58.08 m=2
* device instance $1869 r0 *1 404.54,24.19 dantenna
D$1869 VSS CK4|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1871 r0 *1 504.54,24.19 dantenna
D$1871 VSS CK5|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1873 r0 *1 604.54,24.19 dantenna
D$1873 VSS CK6|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1877 r0 *1 -159.56,320 dantenna
D$1877 VSS IN5|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1878 r0 *1 -159.56,220 dantenna
D$1878 VSS IN6|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1881 r0 *1 -37.46,337.63 dantenna
D$1881 VSS CORE|in5_c dantenna A=1.984 P=7.48 m=1
* device instance $1882 r0 *1 -37.46,237.63 dantenna
D$1882 VSS CORE|in6_c dantenna A=1.984 P=7.48 m=1
* device instance $1883 r0 *1 245.225,142.54 dantenna
D$1883 VSS CORE dantenna A=1.984 P=7.48 m=1
* device instance $1884 r0 *1 445.225,142.54 dantenna
D$1884 VSS CORE$1 dantenna A=1.984 P=7.48 m=1
* device instance $1885 r0 *1 545.225,142.54 dantenna
D$1885 VSS CORE$2 dantenna A=1.984 P=7.48 m=1
* device instance $1886 r0 *1 645.225,142.54 dantenna
D$1886 VSS CORE$3 dantenna A=1.984 P=7.48 m=1
* device instance $1887 r0 *1 935.06,220 dantenna
D$1887 VSS OUT6 dantenna A=35.0028 P=58.08 m=2
* device instance $1888 r0 *1 935.06,320 dantenna
D$1888 VSS OUT5 dantenna A=35.0028 P=58.08 m=2
* device instance $1891 r0 *1 947.17,297.975 dantenna
D$1891 VSS \$357 dantenna A=0.192 P=1.88 m=1
* device instance $1892 r0 *1 947.17,197.975 dantenna
D$1892 VSS \$244 dantenna A=0.192 P=1.88 m=1
* device instance $1893 r0 *1 947.17,397.975 dantenna
D$1893 VSS \$470 dantenna A=0.192 P=1.88 m=1
* device instance $1894 r0 *1 -159.56,420 dantenna
D$1894 VSS IN4|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1896 r0 *1 935.06,420 dantenna
D$1896 VSS OUT4 dantenna A=35.0028 P=58.08 m=2
* device instance $1898 r0 *1 -37.46,437.63 dantenna
D$1898 VSS CORE|in4_c dantenna A=1.984 P=7.48 m=1
* device instance $1901 r0 *1 -159.56,520 dantenna
D$1901 VSS PAD|VLO dantenna A=35.0028 P=58.08 m=2
* device instance $1903 r0 *1 -37.46,537.63 dantenna
D$1903 VSS CORE$4 dantenna A=1.984 P=7.48 m=1
* device instance $1904 r0 *1 932.65,584.765 dantenna
D$1904 VSS \$619 dantenna A=0.192 P=1.88 m=1
* device instance $1905 r0 *1 -159.56,620 dantenna
D$1905 VSS PAD|VHI dantenna A=35.0028 P=58.08 m=2
* device instance $1907 r0 *1 -37.46,637.63 dantenna
D$1907 VSS CORE$5 dantenna A=1.984 P=7.48 m=1
* device instance $1908 r0 *1 947.17,697.975 dantenna
D$1908 VSS \$731 dantenna A=0.192 P=1.88 m=1
* device instance $1909 r0 *1 -159.56,720 dantenna
D$1909 VSS IN3|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1911 r0 *1 935.06,720 dantenna
D$1911 VSS OUT3 dantenna A=35.0028 P=58.08 m=2
* device instance $1913 r0 *1 -37.46,737.63 dantenna
D$1913 VSS CORE|in3_c dantenna A=1.984 P=7.48 m=1
* device instance $1914 r0 *1 947.17,797.975 dantenna
D$1914 VSS \$844 dantenna A=0.192 P=1.88 m=1
* device instance $1915 r0 *1 -159.56,820 dantenna
D$1915 VSS IN2|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1917 r0 *1 935.06,820 dantenna
D$1917 VSS OUT2 dantenna A=35.0028 P=58.08 m=2
* device instance $1919 r0 *1 -37.46,837.63 dantenna
D$1919 VSS CORE|in2_c dantenna A=1.984 P=7.48 m=1
* device instance $1920 r0 *1 947.17,897.975 dantenna
D$1920 VSS \$957 dantenna A=0.192 P=1.88 m=1
* device instance $1921 r0 *1 -159.56,920 dantenna
D$1921 VSS IN1|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1923 r0 *1 935.06,920 dantenna
D$1923 VSS OUT1 dantenna A=35.0028 P=58.08 m=2
* device instance $1925 r0 *1 -37.46,937.63 dantenna
D$1925 VSS CORE|in1_c dantenna A=1.984 P=7.48 m=1
* device instance $1926 r0 *1 157.63,997.46 dantenna
D$1926 VSS CORE|vref_c dantenna A=1.984 P=7.48 m=1
* device instance $1927 r0 *1 257.63,997.46 dantenna
D$1927 VSS CORE$9 dantenna A=1.984 P=7.48 m=1
* device instance $1928 r0 *1 445.225,997.46 dantenna
D$1928 VSS CORE$6 dantenna A=1.984 P=7.48 m=1
* device instance $1929 r0 *1 545.225,997.46 dantenna
D$1929 VSS CORE$7 dantenna A=1.984 P=7.48 m=1
* device instance $1930 r0 *1 645.225,997.46 dantenna
D$1930 VSS CORE$8 dantenna A=1.984 P=7.48 m=1
* device instance $1931 r0 *1 404.54,1115.81 dantenna
D$1931 VSS CK3|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1933 r0 *1 504.54,1115.81 dantenna
D$1933 VSS CK2|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1935 r0 *1 604.54,1115.81 dantenna
D$1935 VSS CK1|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1937 r0 *1 4.765,1112.65 dantenna
D$1937 VSS \$1105 dantenna A=0.192 P=1.88 m=1
* device instance $1938 r0 *1 140,1115.06 dantenna
D$1938 VSS PAD|VREF dantenna A=35.0028 P=58.08 m=2
* device instance $1939 r0 *1 240,1115.06 dantenna
D$1939 VSS PAD|VLDO dantenna A=35.0028 P=58.08 m=2
* device instance $1940 r0 *1 304.765,1112.65 dantenna
D$1940 VSS \$1106 dantenna A=0.192 P=1.88 m=1
* device instance $1941 r0 *1 704.765,1112.65 dantenna
D$1941 VSS \$1107 dantenna A=0.192 P=1.88 m=1
* device instance $1944 r0 *1 4.54,83.19 dpantenna
D$1944 VSS AVDD dpantenna A=35.0028 P=58.08 m=4
* device instance $1948 r0 *1 204.54,83.19 dpantenna
D$1948 PAD|RES IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1950 r0 *1 304.54,83.19 dpantenna
D$1950 VSS IOVDD dpantenna A=35.0028 P=58.08 m=6
* device instance $1952 r0 *1 404.54,83.19 dpantenna
D$1952 CK4|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1954 r0 *1 504.54,83.19 dpantenna
D$1954 CK5|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1956 r0 *1 604.54,83.19 dpantenna
D$1956 CK6|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1960 r0 *1 -32.49,235.46 dpantenna
D$1960 CORE|in6_c AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1961 r0 *1 -32.49,335.46 dpantenna
D$1961 CORE|in5_c AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1962 r0 *1 -32.49,435.46 dpantenna
D$1962 CORE|in4_c AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1963 r0 *1 -32.49,535.46 dpantenna
D$1963 CORE$4 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1964 r0 *1 -32.49,635.46 dpantenna
D$1964 CORE$5 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1965 r0 *1 -32.49,735.46 dpantenna
D$1965 CORE|in3_c AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1966 r0 *1 -32.49,835.46 dpantenna
D$1966 CORE|in2_c AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1967 r0 *1 -32.49,935.46 dpantenna
D$1967 CORE|in1_c AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1968 r0 *1 155.46,992.49 dpantenna
D$1968 CORE|vref_c AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1969 r0 *1 255.46,992.49 dpantenna
D$1969 CORE$9 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1970 r0 *1 243.055,147.51 dpantenna
D$1970 CORE IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1971 r0 *1 443.055,147.51 dpantenna
D$1971 CORE$1 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1972 r0 *1 543.055,147.51 dpantenna
D$1972 CORE$2 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1973 r0 *1 643.055,147.51 dpantenna
D$1973 CORE$3 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1974 r0 *1 443.055,992.49 dpantenna
D$1974 CORE$6 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1975 r0 *1 543.055,992.49 dpantenna
D$1975 CORE$7 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1976 r0 *1 643.055,992.49 dpantenna
D$1976 CORE$8 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1977 r0 *1 878.81,197.975 dpantenna
D$1977 \$208 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $1978 r0 *1 -124.04,220 dpantenna
D$1978 IN6|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1980 r0 *1 899.54,220 dpantenna
D$1980 OUT6 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1982 r0 *1 -124.04,320 dpantenna
D$1982 IN5|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1984 r0 *1 878.81,297.975 dpantenna
D$1984 \$321 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $1985 r0 *1 899.54,320 dpantenna
D$1985 OUT5 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1987 r0 *1 -124.04,420 dpantenna
D$1987 IN4|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1989 r0 *1 878.81,397.975 dpantenna
D$1989 \$434 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $1990 r0 *1 899.54,420 dpantenna
D$1990 OUT4 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1992 r0 *1 -124.04,520 dpantenna
D$1992 PAD|VLO AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1996 r0 *1 -124.04,620 dpantenna
D$1996 PAD|VHI AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1998 r0 *1 878.81,697.975 dpantenna
D$1998 \$695 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $1999 r0 *1 -124.04,720 dpantenna
D$1999 IN3|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2001 r0 *1 899.54,720 dpantenna
D$2001 OUT3 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2003 r0 *1 -124.04,820 dpantenna
D$2003 IN2|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2005 r0 *1 878.81,797.975 dpantenna
D$2005 \$808 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $2006 r0 *1 899.54,820 dpantenna
D$2006 OUT2 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2008 r0 *1 -124.04,920 dpantenna
D$2008 IN1|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2010 r0 *1 878.81,897.975 dpantenna
D$2010 \$921 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $2011 r0 *1 899.54,920 dpantenna
D$2011 OUT1 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2013 r0 *1 404.54,1056.81 dpantenna
D$2013 CK3|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2015 r0 *1 504.54,1056.81 dpantenna
D$2015 CK2|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2017 r0 *1 604.54,1056.81 dpantenna
D$2017 CK1|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2019 r0 *1 140,1079.54 dpantenna
D$2019 PAD|VREF AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2021 r0 *1 240,1079.54 dpantenna
D$2021 PAD|VLDO AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2023 r0 *1 240.685,141.11 rppd
R$2023 PAD|RES CORE rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2024 r0 *1 440.685,141.11 rppd
R$2024 CK4|PAD CORE$1 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2025 r0 *1 540.685,141.11 rppd
R$2025 CK5|PAD CORE$2 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2026 r0 *1 640.685,141.11 rppd
R$2026 CK6|PAD CORE$3 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2027 r0 *1 -171.25,246.305 rppd
R$2027 VSS \$217 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $2028 r0 *1 -112.25,246.305 rppd
R$2028 AVDD \$218 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $2029 r0 *1 -38.89,233.09 rppd
R$2029 IN6|PAD CORE|in6_c rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2030 r0 *1 -171.25,346.305 rppd
R$2030 VSS \$330 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $2031 r0 *1 -112.25,346.305 rppd
R$2031 AVDD \$331 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $2032 r0 *1 -38.89,333.09 rppd
R$2032 IN5|PAD CORE|in5_c rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2033 r0 *1 -171.25,446.305 rppd
R$2033 VSS \$443 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $2034 r0 *1 -112.25,446.305 rppd
R$2034 AVDD \$444 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $2035 r0 *1 -38.89,433.09 rppd
R$2035 IN4|PAD CORE|in4_c rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2036 r0 *1 -171.25,546.305 rppd
R$2036 VSS \$559 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $2037 r0 *1 -112.25,546.305 rppd
R$2037 AVDD \$560 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $2038 r0 *1 -38.89,533.09 rppd
R$2038 PAD|VLO CORE$4 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2039 r0 *1 901.29,598.875 rppd
R$2039 IOVDD \$620 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $2040 r0 *1 -38.89,633.09 rppd
R$2040 PAD|VHI CORE$5 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2041 r0 *1 -171.25,646.305 rppd
R$2041 VSS \$625 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $2042 r0 *1 -112.25,646.305 rppd
R$2042 AVDD \$626 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $2043 r0 *1 -171.25,746.305 rppd
R$2043 VSS \$704 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $2044 r0 *1 -112.25,746.305 rppd
R$2044 AVDD \$705 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $2045 r0 *1 -38.89,733.09 rppd
R$2045 IN3|PAD CORE|in3_c rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2046 r0 *1 -171.25,846.305 rppd
R$2046 VSS \$817 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $2047 r0 *1 -112.25,846.305 rppd
R$2047 AVDD \$818 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $2048 r0 *1 -38.89,833.09 rppd
R$2048 IN2|PAD CORE|in2_c rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2049 r0 *1 -171.25,946.305 rppd
R$2049 VSS \$930 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $2050 r0 *1 -112.25,946.305 rppd
R$2050 AVDD \$931 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $2051 r0 *1 -38.89,933.09 rppd
R$2051 IN1|PAD CORE|in1_c rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2052 r0 *1 153.09,996.03 rppd
R$2052 CORE|vref_c PAD|VREF rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2053 r0 *1 253.09,996.03 rppd
R$2053 CORE$9 PAD|VLDO rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2054 r0 *1 440.685,996.03 rppd
R$2054 CORE$6 CK3|PAD rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2055 r0 *1 540.685,996.03 rppd
R$2055 CORE$7 CK2|PAD rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2056 r0 *1 640.685,996.03 rppd
R$2056 CORE$8 CK1|PAD rppd w=1 l=2 ps=0 b=0 m=1
* device instance $2057 r0 *1 18.875,1081.29 rppd
R$2057 AVDD \$1164 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $2058 r0 *1 166.305,1058.49 rppd
R$2058 \$1122 AVDD rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $2059 r0 *1 266.305,1058.49 rppd
R$2059 \$1123 AVDD rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $2060 r0 *1 318.875,1081.29 rppd
R$2060 IOVDD \$1165 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $2061 r0 *1 718.875,1081.29 rppd
R$2061 VDD \$1166 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $2062 r0 *1 166.305,1126.85 rppd
R$2062 \$1236 VSS rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $2063 r0 *1 266.305,1126.85 rppd
R$2063 \$1237 VSS rppd w=0.5 l=3.54 ps=0 b=0 m=1
.ENDS padring

* Extracted by KLayout with SG13G2 LVS runset on : 28/04/2024 08:25

* cell sg13g2_IOPadAnalog
.SUBCKT sg13g2_IOPadAnalog
* device instance $1 r0 *1 25.52,10.95 sg13_hv_nmos
M$1 vssio vssio PAD vssio sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $2 r0 *1 27.3,10.95 sg13_hv_nmos
M$2 PAD vssio vssio vssio sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $3 r0 *1 28.54,10.95 sg13_hv_nmos
M$3 vssio vssio PAD vssio sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $4 r0 *1 30.32,10.95 sg13_hv_nmos
M$4 PAD vssio vssio vssio sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $5 r0 *1 31.56,10.95 sg13_hv_nmos
M$5 vssio vssio PAD vssio sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $6 r0 *1 33.34,10.95 sg13_hv_nmos
M$6 PAD vssio vssio vssio sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $7 r0 *1 34.58,10.95 sg13_hv_nmos
M$7 vssio vssio PAD vssio sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $8 r0 *1 36.36,10.95 sg13_hv_nmos
M$8 PAD vssio vssio vssio sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $9 r0 *1 37.6,10.95 sg13_hv_nmos
M$9 vssio vssio PAD vssio sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $10 r0 *1 39.38,10.95 sg13_hv_nmos
M$10 PAD vssio vssio vssio sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $11 r0 *1 40.62,10.95 sg13_hv_nmos
M$11 vssio vssio PAD vssio sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $12 r0 *1 42.4,10.95 sg13_hv_nmos
M$12 PAD vssio vssio vssio sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $13 r0 *1 43.64,10.95 sg13_hv_nmos
M$13 vssio vssio PAD vssio sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $14 r0 *1 45.42,10.95 sg13_hv_nmos
M$14 PAD vssio vssio vssio sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $15 r0 *1 46.66,10.95 sg13_hv_nmos
M$15 vssio vssio PAD vssio sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $16 r0 *1 48.44,10.95 sg13_hv_nmos
M$16 PAD vssio vssio vssio sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $17 r0 *1 49.68,10.95 sg13_hv_nmos
M$17 vssio vssio PAD vssio sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $18 r0 *1 51.46,10.95 sg13_hv_nmos
M$18 PAD vssio vssio vssio sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $19 r0 *1 52.7,10.95 sg13_hv_nmos
M$19 vssio vssio PAD vssio sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $20 r0 *1 54.48,10.95 sg13_hv_nmos
M$20 PAD vssio vssio vssio sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $21 r0 *1 25.52,71.08 sg13_hv_pmos
M$21 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $22 r0 *1 27.3,71.08 sg13_hv_pmos
M$22 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $23 r0 *1 28.54,71.08 sg13_hv_pmos
M$23 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $24 r0 *1 30.32,71.08 sg13_hv_pmos
M$24 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $25 r0 *1 31.56,71.08 sg13_hv_pmos
M$25 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $26 r0 *1 33.34,71.08 sg13_hv_pmos
M$26 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $27 r0 *1 34.58,71.08 sg13_hv_pmos
M$27 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $28 r0 *1 36.36,71.08 sg13_hv_pmos
M$28 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $29 r0 *1 37.6,71.08 sg13_hv_pmos
M$29 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $30 r0 *1 39.38,71.08 sg13_hv_pmos
M$30 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $31 r0 *1 40.62,71.08 sg13_hv_pmos
M$31 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $32 r0 *1 42.4,71.08 sg13_hv_pmos
M$32 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $33 r0 *1 43.64,71.08 sg13_hv_pmos
M$33 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $34 r0 *1 45.42,71.08 sg13_hv_pmos
M$34 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $35 r0 *1 46.66,71.08 sg13_hv_pmos
M$35 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $36 r0 *1 48.44,71.08 sg13_hv_pmos
M$36 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $37 r0 *1 49.68,71.08 sg13_hv_pmos
M$37 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $38 r0 *1 51.46,71.08 sg13_hv_pmos
M$38 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $39 r0 *1 52.7,71.08 sg13_hv_pmos
M$39 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $40 r0 *1 54.48,71.08 sg13_hv_pmos
M$40 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $41 r0 *1 25.52,78.18 sg13_hv_pmos
M$41 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $42 r0 *1 27.3,78.18 sg13_hv_pmos
M$42 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $43 r0 *1 28.54,78.18 sg13_hv_pmos
M$43 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $44 r0 *1 30.32,78.18 sg13_hv_pmos
M$44 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $45 r0 *1 31.56,78.18 sg13_hv_pmos
M$45 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $46 r0 *1 33.34,78.18 sg13_hv_pmos
M$46 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $47 r0 *1 34.58,78.18 sg13_hv_pmos
M$47 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $48 r0 *1 36.36,78.18 sg13_hv_pmos
M$48 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $49 r0 *1 37.6,78.18 sg13_hv_pmos
M$49 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $50 r0 *1 39.38,78.18 sg13_hv_pmos
M$50 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $51 r0 *1 40.62,78.18 sg13_hv_pmos
M$51 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $52 r0 *1 42.4,78.18 sg13_hv_pmos
M$52 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $53 r0 *1 43.64,78.18 sg13_hv_pmos
M$53 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $54 r0 *1 45.42,78.18 sg13_hv_pmos
M$54 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $55 r0 *1 46.66,78.18 sg13_hv_pmos
M$55 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $56 r0 *1 48.44,78.18 sg13_hv_pmos
M$56 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $57 r0 *1 49.68,78.18 sg13_hv_pmos
M$57 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $58 r0 *1 51.46,78.18 sg13_hv_pmos
M$58 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $59 r0 *1 52.7,78.18 sg13_hv_pmos
M$59 \$19 \$19 PAD \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $60 r0 *1 54.48,78.18 sg13_hv_pmos
M$60 PAD \$19 \$19 \$19 sg13_hv_pmos W=6.659999999999998 L=0.5999999999999999
* device instance $61 r0 *1 25.52,10.95 rfnmoshv
61$61 vssio vssio PAD vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $62 r0 *1 27.3,10.95 rfnmoshv
62$62 PAD vssio vssio vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $63 r0 *1 28.54,10.95 rfnmoshv
63$63 vssio vssio PAD vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $64 r0 *1 30.32,10.95 rfnmoshv
64$64 PAD vssio vssio vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $65 r0 *1 31.56,10.95 rfnmoshv
65$65 vssio vssio PAD vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $66 r0 *1 33.34,10.95 rfnmoshv
66$66 PAD vssio vssio vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $67 r0 *1 34.58,10.95 rfnmoshv
67$67 vssio vssio PAD vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $68 r0 *1 36.36,10.95 rfnmoshv
68$68 PAD vssio vssio vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $69 r0 *1 37.6,10.95 rfnmoshv
69$69 vssio vssio PAD vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $70 r0 *1 39.38,10.95 rfnmoshv
70$70 PAD vssio vssio vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $71 r0 *1 40.62,10.95 rfnmoshv
71$71 vssio vssio PAD vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $72 r0 *1 42.4,10.95 rfnmoshv
72$72 PAD vssio vssio vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $73 r0 *1 43.64,10.95 rfnmoshv
73$73 vssio vssio PAD vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $74 r0 *1 45.42,10.95 rfnmoshv
74$74 PAD vssio vssio vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $75 r0 *1 46.66,10.95 rfnmoshv
75$75 vssio vssio PAD vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $76 r0 *1 48.44,10.95 rfnmoshv
76$76 PAD vssio vssio vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $77 r0 *1 49.68,10.95 rfnmoshv
77$77 vssio vssio PAD vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $78 r0 *1 51.46,10.95 rfnmoshv
78$78 PAD vssio vssio vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $79 r0 *1 52.7,10.95 rfnmoshv
79$79 vssio vssio PAD vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $80 r0 *1 54.48,10.95 rfnmoshv
80$80 PAD vssio vssio vssio rfnmoshv W=4.3999999999999995 L=0.5999999999999998
* device instance $81 r0 *1 25.52,71.08 rfpmoshv
81$81 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $82 r0 *1 27.3,71.08 rfpmoshv
82$82 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $83 r0 *1 28.54,71.08 rfpmoshv
83$83 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $84 r0 *1 30.32,71.08 rfpmoshv
84$84 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $85 r0 *1 31.56,71.08 rfpmoshv
85$85 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $86 r0 *1 33.34,71.08 rfpmoshv
86$86 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $87 r0 *1 34.58,71.08 rfpmoshv
87$87 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $88 r0 *1 36.36,71.08 rfpmoshv
88$88 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $89 r0 *1 37.6,71.08 rfpmoshv
89$89 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $90 r0 *1 39.38,71.08 rfpmoshv
90$90 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $91 r0 *1 40.62,71.08 rfpmoshv
91$91 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $92 r0 *1 42.4,71.08 rfpmoshv
92$92 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $93 r0 *1 43.64,71.08 rfpmoshv
93$93 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $94 r0 *1 45.42,71.08 rfpmoshv
94$94 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $95 r0 *1 46.66,71.08 rfpmoshv
95$95 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $96 r0 *1 48.44,71.08 rfpmoshv
96$96 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $97 r0 *1 49.68,71.08 rfpmoshv
97$97 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $98 r0 *1 51.46,71.08 rfpmoshv
98$98 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $99 r0 *1 52.7,71.08 rfpmoshv
99$99 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $100 r0 *1 54.48,71.08 rfpmoshv
100$100 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $101 r0 *1 25.52,78.18 rfpmoshv
101$101 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $102 r0 *1 27.3,78.18 rfpmoshv
102$102 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $103 r0 *1 28.54,78.18 rfpmoshv
103$103 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $104 r0 *1 30.32,78.18 rfpmoshv
104$104 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $105 r0 *1 31.56,78.18 rfpmoshv
105$105 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $106 r0 *1 33.34,78.18 rfpmoshv
106$106 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $107 r0 *1 34.58,78.18 rfpmoshv
107$107 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $108 r0 *1 36.36,78.18 rfpmoshv
108$108 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $109 r0 *1 37.6,78.18 rfpmoshv
109$109 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $110 r0 *1 39.38,78.18 rfpmoshv
110$110 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $111 r0 *1 40.62,78.18 rfpmoshv
111$111 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $112 r0 *1 42.4,78.18 rfpmoshv
112$112 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $113 r0 *1 43.64,78.18 rfpmoshv
113$113 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $114 r0 *1 45.42,78.18 rfpmoshv
114$114 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $115 r0 *1 46.66,78.18 rfpmoshv
115$115 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $116 r0 *1 48.44,78.18 rfpmoshv
116$116 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $117 r0 *1 49.68,78.18 rfpmoshv
117$117 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $118 r0 *1 51.46,78.18 rfpmoshv
118$118 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $119 r0 *1 52.7,78.18 rfpmoshv
119$119 \$19 \$19 PAD \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $120 r0 *1 54.48,78.18 rfpmoshv
120$120 PAD \$19 \$19 \$19 rfpmoshv W=6.659999999999998 L=0.5999999999999999
* device instance $121 r0 *1 57.63,142.54 dantenna
D$121 vssio CORE dantenna A=1.984 P=7.48 m=1
* device instance $122 r0 *1 55.46,147.51 dpantenna
D$122 CORE IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $123 r0 *1 53.09,141.11 res_rppd
R$123 PAD CORE res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0 ps=0.0
+ m=1.0
.ENDS sg13g2_IOPadAnalog

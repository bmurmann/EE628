* Extracted by KLayout with SG13G2 LVS runset on : 27/04/2024 01:01

* cell sg13g2_buf_4
.SUBCKT sg13g2_buf_4
* device instance $1 r0 *1 0.62,0.96 sg13_lv_nmos
M$1 sub! \$4 \$3 sub! sg13_lv_nmos W=2.96 L=0.13
* device instance $5 r0 *1 3.1,0.96 sg13_lv_nmos
M$5 sub! \$5 \$4 sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $6 r0 *1 2.66,2.48 sg13_lv_pmos
M$6 \$2 \$5 \$4 \$2 sg13_lv_pmos W=1.68 L=0.13
* device instance $8 r0 *1 0.62,2.62 sg13_lv_pmos
M$8 \$2 \$4 \$3 \$2 sg13_lv_pmos W=4.48 L=0.13
.ENDS sg13g2_buf_4

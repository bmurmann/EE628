* Extracted by KLayout with SG13G2 LVS runset on : 25/05/2024 03:57

* cell UHEE628_S2024
* pin PAD,RES
* pin CK4,PAD
* pin CK5,PAD
* pin CK6,PAD
* pin IOVDD
* pin AVDD
* pin CORE
* pin CORE
* pin CORE
* pin CORE
* pin IN6,PAD
* pin OUT6
* pin VDD
* pin dout
* pin CORE
* pin IN5,PAD
* pin OUT5
* pin CORE
* pin IN4,PAD
* pin OUT4
* pin CORE
* pin PAD,VLO
* pin CORE
* pin PAD,VHI
* pin CORE
* pin IN3,PAD
* pin OUT3
* pin CORE
* pin PAD,VLDO
* pin IN2,PAD
* pin OUT2
* pin CORE
* pin CORE
* pin IN1,PAD
* pin OUT1
* pin CORE
* pin PAD,VREF
* pin CORE
* pin CORE
* pin CORE
* pin CORE
* pin CK3,PAD
* pin CK2,PAD
* pin CK1,PAD
* pin VSS
.SUBCKT UHEE628_S2024 PAD|RES CK4|PAD CK5|PAD CK6|PAD IOVDD AVDD CORE CORE$1
+ CORE$2 CORE$3 IN6|PAD OUT6 VDD dout CORE$4 IN5|PAD OUT5 CORE$5 IN4|PAD OUT4
+ CORE$6 PAD|VLO CORE$7 PAD|VHI CORE$8 IN3|PAD OUT3 CORE$9 PAD|VLDO IN2|PAD
+ OUT2 CORE$10 CORE$11 IN1|PAD OUT1 CORE$12 PAD|VREF CORE$13 CORE$14 CORE$15
+ CORE$16 CK3|PAD CK2|PAD CK1|PAD VSS
* device instance $1 r0 *1 500.255,239.005 sg13_lv_nmos
M$1 \$173 \$178 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $2 r0 *1 700.255,239.005 sg13_lv_nmos
M$2 \$174 \$179 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $3 r0 *1 800.255,239.005 sg13_lv_nmos
M$3 \$175 \$180 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $4 r0 *1 900.255,239.005 sg13_lv_nmos
M$4 \$176 \$181 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $5 r0 *1 1060.995,297.48 sg13_lv_nmos
M$5 \$230 dout VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $6 r0 *1 431.875,301.115 sg13_lv_nmos
M$6 \$261 \$283 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $8 r0 *1 432.905,301.115 sg13_lv_nmos
M$8 \$261 \$374 \$270 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $10 r0 *1 434.755,301.115 sg13_lv_nmos
M$10 \$262 \$284 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $12 r0 *1 435.785,301.115 sg13_lv_nmos
M$12 \$262 \$324 \$263 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $14 r0 *1 437.56,301.14 sg13_lv_nmos
M$14 VSS \$270 \$264 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $18 r0 *1 440.44,301.14 sg13_lv_nmos
M$18 VSS \$263 \$265 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $22 r0 *1 443.26,301.14 sg13_lv_nmos
M$22 VSS \$264 \$266 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $30 r0 *1 448.06,301.14 sg13_lv_nmos
M$30 VSS \$265 \$267 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $38 r0 *1 431.085,305.825 sg13_lv_nmos
M$38 VSS \$176 \$319 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $40 r0 *1 433.06,305.8 sg13_lv_nmos
M$40 \$320 \$319 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $42 r0 *1 434.09,305.8 sg13_lv_nmos
M$42 \$320 \$283 \$331 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $44 r0 *1 435.865,305.825 sg13_lv_nmos
M$44 VSS \$331 \$321 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $48 r0 *1 438.745,305.825 sg13_lv_nmos
M$48 VSS \$321 \$322 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $52 r0 *1 441.625,305.825 sg13_lv_nmos
M$52 VSS \$322 \$323 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $56 r0 *1 444.505,305.825 sg13_lv_nmos
M$56 VSS \$323 \$324 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $60 r0 *1 447.385,305.825 sg13_lv_nmos
M$60 VSS \$324 \$325 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $64 r0 *1 450.265,305.825 sg13_lv_nmos
M$64 VSS \$325 \$284 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $68 r0 *1 456.79,303.21 sg13_lv_nmos
M$68 VSS \$267 \$291 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $69 r0 *1 457.97,303.37 sg13_lv_nmos
M$69 \$294 \$266 \$306 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $70 r0 *1 458.48,303.37 sg13_lv_nmos
M$70 VSS \$247 \$306 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $71 r0 *1 458.99,303.32 sg13_lv_nmos
M$71 VSS \$294 \$295 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $72 r0 *1 460.28,303.305 sg13_lv_nmos
M$72 VSS \$247 \$296 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $73 r0 *1 461.13,303.21 sg13_lv_nmos
M$73 VSS \$266 \$309 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $74 r0 *1 461.44,303.21 sg13_lv_nmos
M$74 \$309 \$296 \$292 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $75 r0 *1 465.4,304.425 sg13_lv_nmos
M$75 \$297 \$325 \$248 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $76 r0 *1 465.91,304.425 sg13_lv_nmos
M$76 \$248 \$266 \$298 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $77 r0 *1 469.22,304.415 sg13_lv_nmos
M$77 \$272 \$267 \$298 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $78 r0 *1 469.73,304.415 sg13_lv_nmos
M$78 \$298 \$173 \$271 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $79 r0 *1 1060.995,300.99 sg13_lv_nmos
M$79 \$268 dout VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $80 r0 *1 431.05,310.475 sg13_lv_nmos
M$80 VSS \$319 \$368 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $82 r0 *1 433.025,310.45 sg13_lv_nmos
M$82 \$369 \$284 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $84 r0 *1 434.055,310.45 sg13_lv_nmos
M$84 \$369 \$368 \$370 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $86 r0 *1 435.83,310.475 sg13_lv_nmos
M$86 VSS \$370 \$371 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $90 r0 *1 438.71,310.475 sg13_lv_nmos
M$90 VSS \$371 \$372 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $94 r0 *1 441.59,310.475 sg13_lv_nmos
M$94 VSS \$372 \$373 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $98 r0 *1 444.47,310.475 sg13_lv_nmos
M$98 VSS \$373 \$374 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $102 r0 *1 447.35,310.475 sg13_lv_nmos
M$102 VSS \$374 \$375 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $106 r0 *1 450.23,310.475 sg13_lv_nmos
M$106 VSS \$375 \$283 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $110 r0 *1 457.825,307.85 sg13_lv_nmos
M$110 \$347 \$295 PAD|VLO VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $111 r0 *1 460.21,307.855 sg13_lv_nmos
M$111 \$347 \$267 \$346 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $112 r0 *1 465.395,308.555 sg13_lv_nmos
M$112 VSS \$297 \$297 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $113 r0 *1 469.615,308.555 sg13_lv_nmos
M$113 VSS \$272 \$271 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $114 r0 *1 431.685,321.635 sg13_lv_nmos
M$114 VSS \$266 \$442 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $115 r0 *1 432.865,321.795 sg13_lv_nmos
M$115 \$446 \$267 \$451 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $116 r0 *1 433.375,321.795 sg13_lv_nmos
M$116 VSS \$439 \$451 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $117 r0 *1 433.885,321.745 sg13_lv_nmos
M$117 VSS \$446 \$443 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $118 r0 *1 435.175,321.73 sg13_lv_nmos
M$118 VSS \$439 \$447 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $119 r0 *1 436.025,321.635 sg13_lv_nmos
M$119 VSS \$267 \$454 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $120 r0 *1 436.335,321.635 sg13_lv_nmos
M$120 \$454 \$447 \$444 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $121 r0 *1 440.295,322.85 sg13_lv_nmos
M$121 \$448 \$375 \$437 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $122 r0 *1 440.805,322.85 sg13_lv_nmos
M$122 \$437 \$267 \$449 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $123 r0 *1 444.115,322.84 sg13_lv_nmos
M$123 \$440 \$266 \$449 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $124 r0 *1 444.625,322.84 sg13_lv_nmos
M$124 \$449 \$173 \$346 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $125 r0 *1 451.1,325.71 sg13_lv_nmos
M$125 VSS \$266 \$467 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $126 r0 *1 452.54,325.71 sg13_lv_nmos
M$126 VSS \$173 \$493 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $127 r0 *1 453.94,325.71 sg13_lv_nmos
M$127 VSS \$494 \$247 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $129 r0 *1 454.96,325.76 sg13_lv_nmos
M$129 VSS \$546 \$494 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $130 r0 *1 456.195,325.53 sg13_lv_nmos
M$130 \$468 \$546 \$475 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $131 r0 *1 456.505,325.53 sg13_lv_nmos
M$131 \$475 \$493 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $132 r0 *1 457.085,325.915 sg13_lv_nmos
M$132 VSS \$495 \$462 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $133 r0 *1 464.925,325.53 sg13_lv_nmos
M$133 \$470 \$471 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $134 r0 *1 465.435,325.53 sg13_lv_nmos
M$134 VSS \$493 \$476 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $135 r0 *1 465.745,325.53 sg13_lv_nmos
M$135 \$476 \$482 \$471 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $136 r0 *1 467.785,325.64 sg13_lv_nmos
M$136 VSS \$482 \$473 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $137 r0 *1 466.765,325.69 sg13_lv_nmos
M$137 VSS \$482 \$472 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $139 r0 *1 468.805,325.69 sg13_lv_nmos
M$139 VSS \$473 \$439 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $141 r0 *1 470.56,325.71 sg13_lv_nmos
M$141 VSS \$439 dout VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $143 r0 *1 432.72,326.275 sg13_lv_nmos
M$143 \$480 \$443 PAD|VLO VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $144 r0 *1 435.105,326.28 sg13_lv_nmos
M$144 \$480 \$266 CORE$4 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $145 r0 *1 440.29,326.98 sg13_lv_nmos
M$145 VSS \$448 \$448 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $146 r0 *1 444.51,326.98 sg13_lv_nmos
M$146 VSS \$440 \$346 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $147 r0 *1 458.175,325.595 sg13_lv_nmos
M$147 VSS \$493 \$479 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $148 r0 *1 458.485,325.595 sg13_lv_nmos
M$148 \$479 \$462 \$469 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $149 r0 *1 459.26,326.32 sg13_lv_nmos
M$149 \$468 \$463 \$495 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $150 r0 *1 459.77,326.32 sg13_lv_nmos
M$150 \$495 \$481 \$469 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $151 r0 *1 460.575,329.87 sg13_lv_nmos
M$151 VSS \$297 \$533 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $152 r0 *1 460.575,330.815 sg13_lv_nmos
M$152 \$533 \$267 \$538 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $153 r0 *1 460.575,331.325 sg13_lv_nmos
M$153 \$538 \$544 \$543 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $154 r0 *1 461.03,325.795 sg13_lv_nmos
M$154 VSS \$463 \$481 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $155 r0 *1 462.13,325.795 sg13_lv_nmos
M$155 VSS \$266 \$463 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $156 r0 *1 463.65,329.87 sg13_lv_nmos
M$156 VSS \$526 \$534 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $157 r0 *1 463.65,330.815 sg13_lv_nmos
M$157 \$534 \$267 \$539 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $158 r0 *1 463.65,331.325 sg13_lv_nmos
M$158 \$539 \$543 \$544 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $159 r0 *1 463.34,325.915 sg13_lv_nmos
M$159 \$482 \$463 \$470 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $160 r0 *1 463.875,325.755 sg13_lv_nmos
M$160 \$462 \$481 \$482 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $161 r0 *1 467.385,330.81 sg13_lv_nmos
M$161 VSS \$544 \$540 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $162 r0 *1 467.385,331.32 sg13_lv_nmos
M$162 \$540 \$546 \$545 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $163 r0 *1 470.52,330.81 sg13_lv_nmos
M$163 VSS \$543 \$541 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $164 r0 *1 470.52,331.32 sg13_lv_nmos
M$164 \$541 \$545 \$546 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $165 r0 *1 457.62,331.325 sg13_lv_nmos
M$165 \$526 \$266 \$271 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $166 r0 *1 464.23,393.71 sg13_lv_nmos
M$166 \$623 \$625 VSS VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $167 r0 *1 464.74,393.76 sg13_lv_nmos
M$167 VSS \$645 \$628 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $168 r0 *1 465.25,393.76 sg13_lv_nmos
M$168 \$628 \$693 \$625 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $169 r0 *1 476.37,393.76 sg13_lv_nmos
M$169 \$626 \$652 \$631 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $170 r0 *1 476.88,393.76 sg13_lv_nmos
M$170 VSS \$627 \$631 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $171 r0 *1 477.39,393.71 sg13_lv_nmos
M$171 VSS \$626 \$624 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $172 r0 *1 459.485,394.65 sg13_lv_nmos
M$172 PAD|VLO \$623 \$632 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $173 r0 *1 482.135,394.65 sg13_lv_nmos
M$173 PAD|VLO \$624 \$659 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $174 r0 *1 1060.995,397.48 sg13_lv_nmos
M$174 \$643 \$645 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $175 r0 *1 458.33,399.375 sg13_lv_nmos
M$175 \$632 \$652 CORE$5 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $176 r0 *1 483.295,399.375 sg13_lv_nmos
M$176 \$799 \$693 \$659 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $177 r0 *1 1060.995,400.99 sg13_lv_nmos
M$177 \$687 \$645 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $178 r0 *1 443.525,403.27 sg13_lv_nmos
M$178 \$754 \$693 \$616 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $179 r0 *1 448.1,403.27 sg13_lv_nmos
M$179 \$616 \$887 \$696 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $180 r0 *1 493.52,403.27 sg13_lv_nmos
M$180 \$697 \$843 \$617 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $181 r0 *1 498.095,403.27 sg13_lv_nmos
M$181 \$617 \$652 \$755 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $182 r0 *1 458.725,405.86 sg13_lv_nmos
M$182 VSS \$652 \$653 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $183 r0 *1 462.07,405.955 sg13_lv_nmos
M$183 VSS \$645 \$721 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $184 r0 *1 462.92,405.86 sg13_lv_nmos
M$184 VSS \$693 \$727 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $185 r0 *1 463.23,405.86 sg13_lv_nmos
M$185 \$727 \$721 \$711 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $186 r0 *1 478.39,405.86 sg13_lv_nmos
M$186 \$712 \$722 \$729 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $187 r0 *1 478.7,405.86 sg13_lv_nmos
M$187 \$729 \$652 VSS VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $188 r0 *1 479.55,405.955 sg13_lv_nmos
M$188 VSS \$627 \$722 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $189 r0 *1 482.9,405.86 sg13_lv_nmos
M$189 \$654 \$693 VSS VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $190 r0 *1 454.04,411.25 sg13_lv_nmos
M$190 \$696 \$696 VSS VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $191 r0 *1 487.58,411.25 sg13_lv_nmos
M$191 VSS \$697 \$697 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $192 r0 *1 454.04,420.795 sg13_lv_nmos
M$192 \$799 \$615 VSS VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $193 r0 *1 487.58,420.795 sg13_lv_nmos
M$193 VSS \$618 \$795 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $194 r0 *1 458.98,423.25 sg13_lv_nmos
M$194 \$799 \$173 \$754 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $195 r0 *1 463.555,423.25 sg13_lv_nmos
M$195 \$754 \$652 \$615 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $196 r0 *1 478.065,423.25 sg13_lv_nmos
M$196 \$618 \$693 \$755 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $197 r0 *1 482.645,423.25 sg13_lv_nmos
M$197 \$755 \$173 \$795 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $198 r0 *1 452.73,430.97 sg13_lv_nmos
M$198 \$838 \$879 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $200 r0 *1 453.76,430.97 sg13_lv_nmos
M$200 \$838 \$888 \$847 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $202 r0 *1 477.92,430.97 sg13_lv_nmos
M$202 \$845 \$844 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $204 r0 *1 478.95,430.97 sg13_lv_nmos
M$204 \$845 \$842 \$848 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $206 r0 *1 455.995,430.995 sg13_lv_nmos
M$206 VSS \$847 \$839 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $210 r0 *1 459.41,430.995 sg13_lv_nmos
M$210 VSS \$839 \$840 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $214 r0 *1 462.645,430.995 sg13_lv_nmos
M$214 VSS \$840 \$841 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $218 r0 *1 466.17,430.995 sg13_lv_nmos
M$218 VSS \$841 \$842 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $222 r0 *1 470.03,430.995 sg13_lv_nmos
M$222 VSS \$842 \$843 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $226 r0 *1 474,430.995 sg13_lv_nmos
M$226 VSS \$843 \$844 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $230 r0 *1 481.6,430.995 sg13_lv_nmos
M$230 VSS \$848 \$846 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $234 r0 *1 485,430.995 sg13_lv_nmos
M$234 VSS \$846 \$693 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $242 r0 *1 446.845,438.965 sg13_lv_nmos
M$242 VSS \$175 \$879 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $244 r0 *1 449.365,438.965 sg13_lv_nmos
M$244 VSS \$879 \$880 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $246 r0 *1 452.01,438.94 sg13_lv_nmos
M$246 \$881 \$880 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $248 r0 *1 453.04,438.94 sg13_lv_nmos
M$248 \$881 \$844 \$882 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $250 r0 *1 455.375,438.965 sg13_lv_nmos
M$250 VSS \$882 \$883 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $254 r0 *1 459.84,438.965 sg13_lv_nmos
M$254 VSS \$883 \$884 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $258 r0 *1 463.255,438.965 sg13_lv_nmos
M$258 VSS \$884 \$885 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $262 r0 *1 466.775,438.965 sg13_lv_nmos
M$262 VSS \$885 \$886 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $266 r0 *1 470.635,438.965 sg13_lv_nmos
M$266 VSS \$886 \$887 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $270 r0 *1 474.605,438.965 sg13_lv_nmos
M$270 VSS \$887 \$888 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $274 r0 *1 478.275,438.94 sg13_lv_nmos
M$274 \$889 \$888 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $276 r0 *1 479.305,438.94 sg13_lv_nmos
M$276 \$889 \$886 \$890 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $278 r0 *1 481.955,438.965 sg13_lv_nmos
M$278 VSS \$890 \$891 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $282 r0 *1 485.355,438.965 sg13_lv_nmos
M$282 VSS \$891 \$652 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $290 r0 *1 450.19,456.17 sg13_lv_nmos
M$290 VSS \$943 \$1041 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $291 r0 *1 450.19,450.37 sg13_lv_nmos
M$291 VSS \$988 \$1010 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $292 r0 *1 449.325,446.44 sg13_lv_nmos
M$292 VSS \$973 \$627 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $294 r0 *1 450.345,446.49 sg13_lv_nmos
M$294 VSS \$1014 \$973 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $295 r0 *1 450.235,453.87 sg13_lv_nmos
M$295 \$1014 \$1044 \$1010 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $296 r0 *1 450.235,459.67 sg13_lv_nmos
M$296 \$1044 \$1014 \$1041 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $297 r0 *1 452.325,446.26 sg13_lv_nmos
M$297 \$953 \$1014 \$963 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $298 r0 *1 452.635,446.26 sg13_lv_nmos
M$298 \$963 \$946 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $299 r0 *1 453.215,446.645 sg13_lv_nmos
M$299 VSS \$974 \$948 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $300 r0 *1 454.305,446.325 sg13_lv_nmos
M$300 VSS \$946 \$964 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $301 r0 *1 454.615,446.325 sg13_lv_nmos
M$301 \$964 \$948 \$954 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $302 r0 *1 455.39,447.05 sg13_lv_nmos
M$302 \$953 \$947 \$974 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $303 r0 *1 455.9,447.05 sg13_lv_nmos
M$303 \$974 \$984 \$954 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $304 r0 *1 457.16,446.525 sg13_lv_nmos
M$304 VSS \$947 \$984 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $305 r0 *1 458.26,446.525 sg13_lv_nmos
M$305 VSS \$652 \$947 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $306 r0 *1 459.47,446.645 sg13_lv_nmos
M$306 \$956 \$947 \$955 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $307 r0 *1 460.005,446.485 sg13_lv_nmos
M$307 \$948 \$984 \$956 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $308 r0 *1 461.055,446.26 sg13_lv_nmos
M$308 \$955 \$957 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $309 r0 *1 461.565,446.26 sg13_lv_nmos
M$309 VSS \$946 \$966 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $310 r0 *1 461.875,446.26 sg13_lv_nmos
M$310 \$966 \$956 \$957 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $311 r0 *1 463.915,446.37 sg13_lv_nmos
M$311 VSS \$956 \$959 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $312 r0 *1 462.895,446.42 sg13_lv_nmos
M$312 VSS \$956 \$958 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $314 r0 *1 464.935,446.42 sg13_lv_nmos
M$314 VSS \$959 \$645 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $316 r0 *1 467.705,446.44 sg13_lv_nmos
M$316 VSS \$173 \$946 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $317 r0 *1 469.14,446.44 sg13_lv_nmos
M$317 VSS \$652 \$960 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $318 r0 *1 469.695,451.055 sg13_lv_nmos
M$318 \$961 \$652 \$795 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $319 r0 *1 479.86,451.33 sg13_lv_nmos
M$319 VSS \$697 \$1003 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $320 r0 *1 479.86,445.67 sg13_lv_nmos
M$320 VSS \$961 \$942 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $321 r0 *1 483.42,453 sg13_lv_nmos
M$321 \$988 \$943 \$1017 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $322 r0 *1 483.42,447.34 sg13_lv_nmos
M$322 \$943 \$988 \$962 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $323 r0 *1 485.065,453 sg13_lv_nmos
M$323 \$1017 \$693 \$1003 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $324 r0 *1 485.065,447.34 sg13_lv_nmos
M$324 \$962 \$693 \$942 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $325 r0 *1 1060.995,497.48 sg13_lv_nmos
M$325 \$1083 \$1085 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $326 r0 *1 1060.995,500.99 sg13_lv_nmos
M$326 \$1111 \$1085 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $327 r0 *1 485.62,504.425 sg13_lv_nmos
M$327 \$1135 \$1145 \$1151 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $328 r0 *1 486.01,504.425 sg13_lv_nmos
M$328 \$1151 \$1136 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $329 r0 *1 486.57,504.425 sg13_lv_nmos
M$329 VSS \$1122 \$1150 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $330 r0 *1 486.925,504.425 sg13_lv_nmos
M$330 \$1150 \$1135 \$1136 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $331 r0 *1 483.98,504.535 sg13_lv_nmos
M$331 VSS \$1133 \$1134 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $332 r0 *1 484.65,504.535 sg13_lv_nmos
M$332 \$1134 \$1128 \$1135 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $333 r0 *1 482.1,504.65 sg13_lv_nmos
M$333 \$1132 \$1145 \$1133 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $334 r0 *1 482.61,504.65 sg13_lv_nmos
M$334 \$1133 \$1128 \$1149 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $335 r0 *1 483,504.65 sg13_lv_nmos
M$335 \$1149 \$1134 \$1148 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $336 r0 *1 483.36,504.65 sg13_lv_nmos
M$336 VSS \$1122 \$1148 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $337 r0 *1 476.77,504.59 sg13_lv_nmos
M$337 VSS \$1305 \$1131 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $338 r0 *1 487.965,504.59 sg13_lv_nmos
M$338 VSS \$1135 \$1137 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $339 r0 *1 489.165,504.495 sg13_lv_nmos
M$339 \$1138 \$1135 VSS VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $340 r0 *1 489.705,504.59 sg13_lv_nmos
M$340 VSS \$1138 \$1139 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $341 r0 *1 491.9,504.59 sg13_lv_nmos
M$341 VSS \$1139 \$1085 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $343 r0 *1 494.695,504.59 sg13_lv_nmos
M$343 VSS \$173 \$1122 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $344 r0 *1 496.61,504.59 sg13_lv_nmos
M$344 VSS \$1152 \$1140 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $346 r0 *1 497.63,504.64 sg13_lv_nmos
M$346 VSS \$1204 \$1152 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $347 r0 *1 478.82,504.45 sg13_lv_nmos
M$347 \$1132 \$1204 \$1147 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $348 r0 *1 479.19,504.45 sg13_lv_nmos
M$348 \$1147 \$1122 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $349 r0 *1 480.335,504.765 sg13_lv_nmos
M$349 VSS \$1305 \$1145 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $350 r0 *1 480.845,504.765 sg13_lv_nmos
M$350 VSS \$1145 \$1128 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $351 r0 *1 481.505,510.995 sg13_lv_nmos
M$351 VSS \$1189 \$1192 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $352 r0 *1 481.705,513.1 sg13_lv_nmos
M$352 \$1192 \$1243 \$1198 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $353 r0 *1 483.505,509.465 sg13_lv_nmos
M$353 \$1182 \$1305 \$1183 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $354 r0 *1 482.905,513.1 sg13_lv_nmos
M$354 \$1198 \$1200 \$1199 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $355 r0 *1 484.105,513.1 sg13_lv_nmos
M$355 \$1200 \$1199 \$1201 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $356 r0 *1 485.505,510.995 sg13_lv_nmos
M$356 VSS \$1183 \$1193 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $357 r0 *1 485.305,513.1 sg13_lv_nmos
M$357 \$1201 \$1243 \$1193 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $358 r0 *1 488.56,513.1 sg13_lv_nmos
M$358 VSS \$1200 \$1202 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $359 r0 *1 489.76,513.1 sg13_lv_nmos
M$359 \$1202 \$1204 \$1203 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $360 r0 *1 490.96,513.1 sg13_lv_nmos
M$360 \$1204 \$1203 \$1205 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $361 r0 *1 492.16,513.1 sg13_lv_nmos
M$361 \$1205 \$1199 VSS VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $362 r0 *1 438.155,518.845 sg13_lv_nmos
M$362 VSS \$1234 \$1235 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $366 r0 *1 441.035,518.845 sg13_lv_nmos
M$366 VSS \$1235 \$1236 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $370 r0 *1 443.915,518.845 sg13_lv_nmos
M$370 VSS \$1236 \$1237 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $374 r0 *1 446.795,518.845 sg13_lv_nmos
M$374 VSS \$1237 \$1238 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $378 r0 *1 449.675,518.845 sg13_lv_nmos
M$378 VSS \$1238 \$1239 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $382 r0 *1 452.555,518.845 sg13_lv_nmos
M$382 VSS \$1239 \$1240 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $386 r0 *1 458.315,518.845 sg13_lv_nmos
M$386 VSS \$1241 \$1242 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $390 r0 *1 461.135,518.845 sg13_lv_nmos
M$390 VSS \$1242 \$1243 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $398 r0 *1 431.455,521.28 sg13_lv_nmos
M$398 VSS \$174 \$1249 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $400 r0 *1 433.375,521.28 sg13_lv_nmos
M$400 VSS \$1249 \$1295 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $402 r0 *1 435.35,521.255 sg13_lv_nmos
M$402 \$1296 \$1240 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $404 r0 *1 436.38,521.255 sg13_lv_nmos
M$404 \$1296 \$1295 \$1308 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $406 r0 *1 435.35,518.87 sg13_lv_nmos
M$406 \$1264 \$1302 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $408 r0 *1 436.38,518.87 sg13_lv_nmos
M$408 \$1264 \$1249 \$1234 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $410 r0 *1 438.155,521.28 sg13_lv_nmos
M$410 VSS \$1308 \$1297 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $414 r0 *1 441.035,521.28 sg13_lv_nmos
M$414 VSS \$1297 \$1298 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $418 r0 *1 443.915,521.28 sg13_lv_nmos
M$418 VSS \$1298 \$1299 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $422 r0 *1 446.795,521.28 sg13_lv_nmos
M$422 VSS \$1299 \$1300 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $426 r0 *1 449.675,521.28 sg13_lv_nmos
M$426 VSS \$1300 \$1301 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $430 r0 *1 452.555,521.28 sg13_lv_nmos
M$430 VSS \$1301 \$1302 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $434 r0 *1 455.51,518.87 sg13_lv_nmos
M$434 \$1265 \$1240 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $436 r0 *1 456.54,518.87 sg13_lv_nmos
M$436 \$1265 \$1238 \$1241 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $438 r0 *1 455.51,521.255 sg13_lv_nmos
M$438 \$1303 \$1302 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $440 r0 *1 456.54,521.255 sg13_lv_nmos
M$440 \$1303 \$1300 \$1309 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $442 r0 *1 458.315,521.28 sg13_lv_nmos
M$442 VSS \$1309 \$1304 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $446 r0 *1 461.135,521.28 sg13_lv_nmos
M$446 VSS \$1304 \$1305 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $454 r0 *1 431.5,535.26 sg13_lv_nmos
M$454 VSS \$1305 \$1351 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $455 r0 *1 432.935,535.355 sg13_lv_nmos
M$455 VSS \$1139 \$1352 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $456 r0 *1 433.785,535.26 sg13_lv_nmos
M$456 VSS \$1243 \$1370 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $457 r0 *1 434.095,535.26 sg13_lv_nmos
M$457 \$1370 \$1352 \$1353 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $458 r0 *1 434.07,553.205 sg13_lv_nmos
M$458 \$1401 \$1355 PAD|VLO VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $459 r0 *1 435.785,535.42 sg13_lv_nmos
M$459 \$1354 \$1243 \$1368 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $460 r0 *1 436.295,535.42 sg13_lv_nmos
M$460 VSS \$1139 \$1368 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $461 r0 *1 436.805,535.37 sg13_lv_nmos
M$461 VSS \$1354 \$1355 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $462 r0 *1 436.815,553.215 sg13_lv_nmos
M$462 \$1401 \$1305 CORE$6 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $463 r0 *1 443.55,535.275 sg13_lv_nmos
M$463 VSS \$1356 \$1356 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $464 r0 *1 444.09,553.17 sg13_lv_nmos
M$464 \$1356 \$1301 \$1412 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $465 r0 *1 449.83,597.155 sg13_lv_nmos
M$465 \$1478 \$1532 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $467 r0 *1 450.86,597.155 sg13_lv_nmos
M$467 \$1478 \$1488 \$1489 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $469 r0 *1 455.2,535.26 sg13_lv_nmos
M$469 VSS \$1377 \$1372 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $470 r0 *1 454.14,553.165 sg13_lv_nmos
M$470 \$1412 \$1243 \$1414 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $471 r0 *1 455.45,553.165 sg13_lv_nmos
M$471 \$1414 \$1305 \$1377 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $472 r0 *1 456.765,553.165 sg13_lv_nmos
M$472 \$1414 \$173 \$1372 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $473 r0 *1 466.5,535.26 sg13_lv_nmos
M$473 VSS \$1243 \$1357 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $474 r0 *1 467.935,535.355 sg13_lv_nmos
M$474 VSS \$1140 \$1358 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $475 r0 *1 468.785,535.26 sg13_lv_nmos
M$475 VSS \$1305 \$1365 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $476 r0 *1 469.095,535.26 sg13_lv_nmos
M$476 \$1365 \$1358 \$1359 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $477 r0 *1 469.07,553.205 sg13_lv_nmos
M$477 \$1402 \$1361 PAD|VLO VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $478 r0 *1 469.99,597.155 sg13_lv_nmos
M$478 \$1485 \$1484 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $480 r0 *1 471.02,597.155 sg13_lv_nmos
M$480 \$1485 \$1482 \$1490 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $482 r0 *1 470.785,535.42 sg13_lv_nmos
M$482 \$1360 \$1305 \$1363 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $483 r0 *1 471.295,535.42 sg13_lv_nmos
M$483 VSS \$1140 \$1363 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $484 r0 *1 471.805,535.37 sg13_lv_nmos
M$484 VSS \$1360 \$1361 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $485 r0 *1 471.815,553.215 sg13_lv_nmos
M$485 \$1402 \$1243 \$1372 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $486 r0 *1 478.55,535.275 sg13_lv_nmos
M$486 VSS \$1189 \$1189 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $487 r0 *1 479.09,553.17 sg13_lv_nmos
M$487 \$1189 \$1239 \$1413 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $488 r0 *1 490.2,535.26 sg13_lv_nmos
M$488 VSS \$1378 \$1182 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $489 r0 *1 489.14,553.165 sg13_lv_nmos
M$489 \$1413 \$1305 \$1411 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $490 r0 *1 490.45,553.165 sg13_lv_nmos
M$490 \$1411 \$1243 \$1378 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $491 r0 *1 491.765,553.165 sg13_lv_nmos
M$491 \$1411 \$173 \$1182 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $492 r0 *1 452.635,597.18 sg13_lv_nmos
M$492 VSS \$1489 \$1479 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $496 r0 *1 455.515,597.18 sg13_lv_nmos
M$496 VSS \$1479 \$1480 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $500 r0 *1 458.395,597.18 sg13_lv_nmos
M$500 VSS \$1480 \$1481 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $504 r0 *1 461.275,597.18 sg13_lv_nmos
M$504 VSS \$1481 \$1482 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $508 r0 *1 464.155,597.18 sg13_lv_nmos
M$508 VSS \$1482 \$1483 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $512 r0 *1 467.035,597.18 sg13_lv_nmos
M$512 VSS \$1483 \$1484 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $516 r0 *1 472.795,597.18 sg13_lv_nmos
M$516 VSS \$1490 \$1486 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $520 r0 *1 475.615,597.18 sg13_lv_nmos
M$520 VSS \$1486 \$1487 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $528 r0 *1 445.935,602.98 sg13_lv_nmos
M$528 VSS \$1474 \$1488 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $530 r0 *1 447.855,602.98 sg13_lv_nmos
M$530 VSS \$1488 \$1524 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $532 r0 *1 449.83,602.955 sg13_lv_nmos
M$532 \$1525 \$1484 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $534 r0 *1 450.86,602.955 sg13_lv_nmos
M$534 \$1525 \$1524 \$1526 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $536 r0 *1 452.635,602.98 sg13_lv_nmos
M$536 VSS \$1526 \$1527 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $540 r0 *1 455.515,602.98 sg13_lv_nmos
M$540 VSS \$1527 \$1528 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $544 r0 *1 458.395,602.98 sg13_lv_nmos
M$544 VSS \$1528 \$1529 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $548 r0 *1 461.275,602.98 sg13_lv_nmos
M$548 VSS \$1529 \$1530 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $552 r0 *1 464.155,602.98 sg13_lv_nmos
M$552 VSS \$1530 \$1531 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $556 r0 *1 467.035,602.98 sg13_lv_nmos
M$556 VSS \$1531 \$1532 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $560 r0 *1 469.99,602.955 sg13_lv_nmos
M$560 \$1533 \$1532 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $562 r0 *1 471.02,602.955 sg13_lv_nmos
M$562 \$1533 \$1530 \$1534 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $564 r0 *1 472.795,602.98 sg13_lv_nmos
M$564 VSS \$1534 \$1535 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $568 r0 *1 475.615,602.98 sg13_lv_nmos
M$568 VSS \$1535 \$1536 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $576 r0 *1 433.27,616.415 sg13_lv_nmos
M$576 VSS \$1536 \$1594 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $577 r0 *1 434.36,616.51 sg13_lv_nmos
M$577 VSS \$1567 \$1598 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $578 r0 *1 435.21,616.415 sg13_lv_nmos
M$578 VSS \$1487 \$1607 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $579 r0 *1 435.52,616.415 sg13_lv_nmos
M$579 \$1607 \$1598 \$1595 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $580 r0 *1 436.85,616.575 sg13_lv_nmos
M$580 \$1603 \$1487 \$1615 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $581 r0 *1 437.36,616.575 sg13_lv_nmos
M$581 VSS \$1567 \$1615 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $582 r0 *1 437.87,616.525 sg13_lv_nmos
M$582 VSS \$1603 \$1587 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $583 r0 *1 441.655,618.475 sg13_lv_nmos
M$583 PAD|VLO \$1587 \$1653 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $584 r0 *1 454.37,617.83 sg13_lv_nmos
M$584 \$1723 \$1536 \$1689 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $585 r0 *1 454.37,618.34 sg13_lv_nmos
M$585 \$1689 \$173 \$1633 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $586 r0 *1 454.37,616.04 sg13_lv_nmos
M$586 \$1588 \$1531 \$1612 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $587 r0 *1 454.37,616.55 sg13_lv_nmos
M$587 \$1612 \$1487 \$1689 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $588 r0 *1 469.325,616.415 sg13_lv_nmos
M$588 VSS \$1487 \$1596 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $589 r0 *1 470.415,616.51 sg13_lv_nmos
M$589 VSS \$1568 \$1599 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $590 r0 *1 471.265,616.415 sg13_lv_nmos
M$590 VSS \$1536 \$1610 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $591 r0 *1 471.575,616.415 sg13_lv_nmos
M$591 \$1610 \$1599 \$1597 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $592 r0 *1 472.905,616.575 sg13_lv_nmos
M$592 \$1604 \$1536 \$1622 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $593 r0 *1 473.415,616.575 sg13_lv_nmos
M$593 VSS \$1568 \$1622 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $594 r0 *1 473.925,616.525 sg13_lv_nmos
M$594 VSS \$1604 \$1589 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $595 r0 *1 477.71,618.475 sg13_lv_nmos
M$595 PAD|VLO \$1589 \$1654 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $596 r0 *1 490.425,617.83 sg13_lv_nmos
M$596 \$1724 \$1487 \$1690 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $597 r0 *1 490.425,618.34 sg13_lv_nmos
M$597 \$1690 \$173 \$1634 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $598 r0 *1 490.425,616.04 sg13_lv_nmos
M$598 \$1590 \$1483 \$1613 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $599 r0 *1 490.425,616.55 sg13_lv_nmos
M$599 \$1613 \$1536 \$1690 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $600 r0 *1 505.425,616.53 sg13_lv_nmos
M$600 VSS \$1536 \$1600 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $601 r0 *1 520.915,619.83 sg13_lv_nmos
M$601 \$1665 \$1664 \$1667 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $602 r0 *1 521.225,619.83 sg13_lv_nmos
M$602 \$1667 \$1649 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $603 r0 *1 521.805,620.215 sg13_lv_nmos
M$603 VSS \$1680 \$1655 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $604 r0 *1 522.895,619.895 sg13_lv_nmos
M$604 VSS \$1649 \$1668 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $605 r0 *1 523.205,619.895 sg13_lv_nmos
M$605 \$1668 \$1655 \$1663 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $606 r0 *1 528.06,620.215 sg13_lv_nmos
M$606 \$1666 \$1656 \$1657 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $607 r0 *1 528.595,620.055 sg13_lv_nmos
M$607 \$1655 \$1691 \$1666 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $608 r0 *1 529.645,619.83 sg13_lv_nmos
M$608 \$1657 \$1658 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $609 r0 *1 530.155,619.83 sg13_lv_nmos
M$609 VSS \$1649 \$1670 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $610 r0 *1 530.465,619.83 sg13_lv_nmos
M$610 \$1670 \$1666 \$1658 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $611 r0 *1 532.505,619.94 sg13_lv_nmos
M$611 VSS \$1666 \$1660 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $612 r0 *1 531.485,619.99 sg13_lv_nmos
M$612 VSS \$1666 \$1659 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $614 r0 *1 533.525,619.99 sg13_lv_nmos
M$614 VSS \$1660 \$1567 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $616 r0 *1 535.21,620.01 sg13_lv_nmos
M$616 VSS \$1567 \$1911 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $618 r0 *1 537,620.01 sg13_lv_nmos
M$618 \$1649 \$173 VSS VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $619 r0 *1 433.495,621.675 sg13_lv_nmos
M$619 CORE$9 \$1536 \$1653 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $620 r0 *1 456.64,623.065 sg13_lv_nmos
M$620 VSS \$1723 \$1633 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $621 r0 *1 462.64,623.065 sg13_lv_nmos
M$621 VSS \$1588 \$1588 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $622 r0 *1 469.55,621.675 sg13_lv_nmos
M$622 \$1633 \$1487 \$1654 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $623 r0 *1 492.695,623.065 sg13_lv_nmos
M$623 VSS \$1724 \$1634 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $624 r0 *1 498.695,623.065 sg13_lv_nmos
M$624 VSS \$1590 \$1590 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $625 r0 *1 505.05,623.5 sg13_lv_nmos
M$625 \$1679 \$1536 \$1634 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $626 r0 *1 509.96,626.51 sg13_lv_nmos
M$626 VSS \$1590 \$1731 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $627 r0 *1 514.885,626.51 sg13_lv_nmos
M$627 VSS \$1679 \$1732 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $628 r0 *1 523.98,620.62 sg13_lv_nmos
M$628 \$1665 \$1656 \$1680 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $629 r0 *1 524.49,620.62 sg13_lv_nmos
M$629 \$1680 \$1691 \$1663 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $630 r0 *1 525.75,620.095 sg13_lv_nmos
M$630 VSS \$1656 \$1691 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $631 r0 *1 526.85,620.095 sg13_lv_nmos
M$631 VSS \$1536 \$1656 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $632 r0 *1 532.795,625.47 sg13_lv_nmos
M$632 VSS \$1721 \$1568 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $634 r0 *1 532.845,626.49 sg13_lv_nmos
M$634 VSS \$1664 \$1721 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $635 r0 *1 522.75,627.29 sg13_lv_nmos
M$635 VSS \$1752 \$1737 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $636 r0 *1 529.69,627.28 sg13_lv_nmos
M$636 VSS \$1751 \$1738 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $637 r0 *1 509.855,627.99 sg13_lv_nmos
M$637 \$1731 \$1487 \$1741 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $638 r0 *1 514.795,627.99 sg13_lv_nmos
M$638 \$1732 \$1487 \$1742 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $639 r0 *1 523.03,628.795 sg13_lv_nmos
M$639 \$1737 \$1664 \$1747 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $640 r0 *1 529.34,628.76 sg13_lv_nmos
M$640 \$1738 \$1747 \$1664 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $641 r0 *1 509.835,629.77 sg13_lv_nmos
M$641 \$1741 \$1752 \$1751 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $642 r0 *1 514.62,629.77 sg13_lv_nmos
M$642 \$1742 \$1751 \$1752 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $643 r0 *1 1060.995,797.48 sg13_lv_nmos
M$643 \$1909 \$1911 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $644 r0 *1 1060.995,800.99 sg13_lv_nmos
M$644 \$1937 \$1911 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $645 r0 *1 633.21,835.705 sg13_lv_nmos
M$645 VSS \$2141 \$2141 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $647 r0 *1 630.06,842.755 sg13_lv_nmos
M$647 \$2209 \$2281 \$2174 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $649 r0 *1 622.76,843.455 sg13_lv_nmos
M$649 VSS \$2141 \$2216 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $651 r0 *1 626.34,843.455 sg13_lv_nmos
M$651 VSS \$2174 \$2217 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $653 r0 *1 623.505,845.055 sg13_lv_nmos
M$653 \$2216 \$2339 \$2232 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $655 r0 *1 626.465,845.055 sg13_lv_nmos
M$655 \$2217 \$2339 \$2233 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $657 r0 *1 632.73,845.055 sg13_lv_nmos
M$657 VSS \$2247 \$2234 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $659 r0 *1 635.69,845.055 sg13_lv_nmos
M$659 VSS \$2248 \$2235 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $661 r0 *1 592.87,846.075 sg13_lv_nmos
M$661 VSS \$2180 \$2164 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $663 r0 *1 614.46,846.075 sg13_lv_nmos
M$663 VSS \$2181 \$2209 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $665 r0 *1 623.505,846.655 sg13_lv_nmos
M$665 \$2232 \$2247 \$2248 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $667 r0 *1 626.465,846.655 sg13_lv_nmos
M$667 \$2233 \$2248 \$2247 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $669 r0 *1 632.73,846.655 sg13_lv_nmos
M$669 \$2234 \$2249 \$2258 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $671 r0 *1 635.69,846.655 sg13_lv_nmos
M$671 \$2235 \$2258 \$2249 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $673 r0 *1 585.345,846.75 sg13_lv_nmos
M$673 \$2256 \$2281 CORE$11 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $675 r0 *1 586.14,851.955 sg13_lv_nmos
M$675 PAD|VLO \$2394 \$2256 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $676 r0 *1 588.475,849.385 sg13_lv_nmos
M$676 \$2172 \$2339 \$2261 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $677 r0 *1 588.475,852.475 sg13_lv_nmos
M$677 \$2172 \$2281 \$2180 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $678 r0 *1 589.55,849.385 sg13_lv_nmos
M$678 \$2261 \$2647 \$2141 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $679 r0 *1 606.935,846.735 sg13_lv_nmos
M$679 \$2257 \$2339 \$2164 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $681 r0 *1 607.73,851.955 sg13_lv_nmos
M$681 PAD|VLO \$2395 \$2257 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $682 r0 *1 610.065,852.475 sg13_lv_nmos
M$682 \$2173 \$2339 \$2181 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $683 r0 *1 610.065,849.385 sg13_lv_nmos
M$683 \$2173 \$2281 \$2262 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $684 r0 *1 611.14,849.385 sg13_lv_nmos
M$684 \$2262 \$2314 \$2141 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $685 r0 *1 623.635,852.165 sg13_lv_nmos
M$685 \$2386 \$2249 \$2446 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $686 r0 *1 623.945,852.165 sg13_lv_nmos
M$686 \$2446 \$2385 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $687 r0 *1 624.525,852.55 sg13_lv_nmos
M$687 VSS \$2458 \$2340 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $688 r0 *1 632.365,852.165 sg13_lv_nmos
M$688 \$2387 \$2388 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $689 r0 *1 632.875,852.165 sg13_lv_nmos
M$689 VSS \$2385 \$2450 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $690 r0 *1 633.185,852.165 sg13_lv_nmos
M$690 \$2450 \$2398 \$2388 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $691 r0 *1 635.225,852.275 sg13_lv_nmos
M$691 VSS \$2398 \$2390 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $692 r0 *1 634.205,852.325 sg13_lv_nmos
M$692 VSS \$2398 \$2389 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $694 r0 *1 636.245,852.325 sg13_lv_nmos
M$694 VSS \$2390 \$2561 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $696 r0 *1 620.94,852.345 sg13_lv_nmos
M$696 VSS \$2281 \$2263 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $697 r0 *1 622.38,852.345 sg13_lv_nmos
M$697 VSS \$173 \$2385 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $698 r0 *1 625.615,852.23 sg13_lv_nmos
M$698 VSS \$2385 \$2447 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $699 r0 *1 625.925,852.23 sg13_lv_nmos
M$699 \$2447 \$2340 \$2396 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $700 r0 *1 626.7,852.955 sg13_lv_nmos
M$700 \$2386 \$2341 \$2458 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $701 r0 *1 627.21,852.955 sg13_lv_nmos
M$701 \$2458 \$2397 \$2396 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $702 r0 *1 628.47,852.43 sg13_lv_nmos
M$702 VSS \$2341 \$2397 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $703 r0 *1 629.57,852.43 sg13_lv_nmos
M$703 VSS \$2281 \$2341 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $704 r0 *1 630.78,852.55 sg13_lv_nmos
M$704 \$2398 \$2341 \$2387 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $705 r0 *1 631.315,852.39 sg13_lv_nmos
M$705 \$2340 \$2397 \$2398 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $706 r0 *1 637.86,852.395 sg13_lv_nmos
M$706 VSS \$2249 \$2399 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $707 r0 *1 638.37,852.345 sg13_lv_nmos
M$707 VSS \$2399 \$2562 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $709 r0 *1 640.4,852.345 sg13_lv_nmos
M$709 VSS \$2561 \$2391 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $711 r0 *1 594.145,854.805 sg13_lv_nmos
M$711 \$2172 \$173 \$2164 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $715 r0 *1 615.735,854.805 sg13_lv_nmos
M$715 \$2173 \$173 \$2209 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $719 r0 *1 617.465,863.425 sg13_lv_nmos
M$719 \$2563 \$2597 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $721 r0 *1 618.495,863.425 sg13_lv_nmos
M$721 \$2563 \$2598 \$2578 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $723 r0 *1 640.7,863.425 sg13_lv_nmos
M$723 \$2569 \$2568 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $725 r0 *1 641.73,863.425 sg13_lv_nmos
M$725 \$2569 \$2567 \$2579 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $727 r0 *1 620.495,863.45 sg13_lv_nmos
M$727 VSS \$2578 \$2564 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $731 r0 *1 623.375,863.45 sg13_lv_nmos
M$731 VSS \$2564 \$2565 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $735 r0 *1 626.255,863.45 sg13_lv_nmos
M$735 VSS \$2565 \$2566 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $739 r0 *1 629.135,863.45 sg13_lv_nmos
M$739 VSS \$2566 \$2567 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $743 r0 *1 632.715,863.45 sg13_lv_nmos
M$743 VSS \$2567 \$2314 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $747 r0 *1 636.295,863.45 sg13_lv_nmos
M$747 VSS \$2314 \$2568 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $751 r0 *1 643.75,863.45 sg13_lv_nmos
M$751 VSS \$2579 \$2570 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $755 r0 *1 646.57,863.45 sg13_lv_nmos
M$755 VSS \$2570 \$2339 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $763 r0 *1 577.495,864.355 sg13_lv_nmos
M$763 \$2593 \$2339 \$2607 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $764 r0 *1 578.005,864.355 sg13_lv_nmos
M$764 VSS \$2561 \$2607 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $765 r0 *1 578.515,864.305 sg13_lv_nmos
M$765 VSS \$2593 \$2394 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $766 r0 *1 579.805,864.29 sg13_lv_nmos
M$766 VSS \$2561 \$2594 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $767 r0 *1 580.655,864.195 sg13_lv_nmos
M$767 VSS \$2339 \$2600 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $768 r0 *1 580.965,864.195 sg13_lv_nmos
M$768 \$2600 \$2594 \$2456 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $769 r0 *1 582.555,864.195 sg13_lv_nmos
M$769 VSS \$2281 \$2335 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $770 r0 *1 599.085,864.355 sg13_lv_nmos
M$770 \$2595 \$2281 \$2606 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $771 r0 *1 599.595,864.355 sg13_lv_nmos
M$771 VSS \$2562 \$2606 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $772 r0 *1 600.105,864.305 sg13_lv_nmos
M$772 VSS \$2595 \$2395 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $773 r0 *1 601.395,864.29 sg13_lv_nmos
M$773 VSS \$2562 \$2596 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $774 r0 *1 602.245,864.195 sg13_lv_nmos
M$774 VSS \$2281 \$2603 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $775 r0 *1 602.555,864.195 sg13_lv_nmos
M$775 \$2603 \$2596 \$2457 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $776 r0 *1 604.145,864.195 sg13_lv_nmos
M$776 VSS \$2339 \$2336 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $777 r0 *1 613.57,869.125 sg13_lv_nmos
M$777 VSS \$2651 \$2598 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $779 r0 *1 615.49,869.125 sg13_lv_nmos
M$779 VSS \$2598 \$2640 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $781 r0 *1 617.465,869.1 sg13_lv_nmos
M$781 \$2641 \$2568 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $783 r0 *1 618.495,869.1 sg13_lv_nmos
M$783 \$2641 \$2640 \$2642 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $785 r0 *1 620.495,869.125 sg13_lv_nmos
M$785 VSS \$2642 \$2643 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $789 r0 *1 623.375,869.125 sg13_lv_nmos
M$789 VSS \$2643 \$2644 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $793 r0 *1 626.255,869.125 sg13_lv_nmos
M$793 VSS \$2644 \$2645 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $797 r0 *1 629.135,869.125 sg13_lv_nmos
M$797 VSS \$2645 \$2646 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $801 r0 *1 632.715,869.125 sg13_lv_nmos
M$801 VSS \$2646 \$2647 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $805 r0 *1 636.295,869.125 sg13_lv_nmos
M$805 VSS \$2647 \$2597 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $809 r0 *1 640.44,869.1 sg13_lv_nmos
M$809 \$2648 \$2597 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $811 r0 *1 641.47,869.1 sg13_lv_nmos
M$811 \$2648 \$2646 \$2649 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $813 r0 *1 643.505,869.125 sg13_lv_nmos
M$813 VSS \$2649 \$2650 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $817 r0 *1 646.325,869.125 sg13_lv_nmos
M$817 VSS \$2650 \$2281 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $825 r0 *1 478.38,941.225 sg13_lv_nmos
M$825 VSS \$3100 \$2883 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $826 r0 *1 478.38,936.465 sg13_lv_nmos
M$826 \$2861 \$2863 \$3050 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $827 r0 *1 480.98,941.225 sg13_lv_nmos
M$827 VSS \$2861 \$2884 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $828 r0 *1 483.425,932.84 sg13_lv_nmos
M$828 VSS \$2863 \$2859 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $829 r0 *1 488.24,942.64 sg13_lv_nmos
M$829 VSS \$2942 \$2900 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $830 r0 *1 491.05,942.61 sg13_lv_nmos
M$830 VSS \$2943 \$2901 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $831 r0 *1 503.35,942.605 sg13_lv_nmos
M$831 VSS \$173 \$2885 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $832 r0 *1 504.605,942.425 sg13_lv_nmos
M$832 \$2892 \$2932 \$2920 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $833 r0 *1 504.915,942.425 sg13_lv_nmos
M$833 \$2920 \$2885 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $834 r0 *1 505.495,942.81 sg13_lv_nmos
M$834 VSS \$2935 \$2886 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $835 r0 *1 506.585,942.49 sg13_lv_nmos
M$835 VSS \$2885 \$2922 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $836 r0 *1 506.895,942.49 sg13_lv_nmos
M$836 \$2922 \$2886 \$2902 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $837 r0 *1 509.44,942.69 sg13_lv_nmos
M$837 VSS \$2887 \$2903 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $838 r0 *1 510.54,942.69 sg13_lv_nmos
M$838 VSS \$2863 \$2887 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $839 r0 *1 511.75,942.81 sg13_lv_nmos
M$839 \$2904 \$2887 \$2893 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $840 r0 *1 512.285,942.65 sg13_lv_nmos
M$840 \$2886 \$2903 \$2904 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $841 r0 *1 513.335,942.425 sg13_lv_nmos
M$841 \$2893 \$2894 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $842 r0 *1 513.845,942.425 sg13_lv_nmos
M$842 VSS \$2885 \$2927 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $843 r0 *1 514.155,942.425 sg13_lv_nmos
M$843 \$2927 \$2904 \$2894 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $844 r0 *1 516.195,942.535 sg13_lv_nmos
M$844 VSS \$2904 \$2896 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $845 r0 *1 515.175,942.585 sg13_lv_nmos
M$845 VSS \$2904 \$2895 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $847 r0 *1 517.215,942.585 sg13_lv_nmos
M$847 VSS \$2896 \$2897 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $849 r0 *1 1060.995,900.99 sg13_lv_nmos
M$849 \$2800 \$2391 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $850 r0 *1 1060.995,897.48 sg13_lv_nmos
M$850 \$2773 \$2391 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $851 r0 *1 441.615,944.16 sg13_lv_nmos
M$851 VSS \$2873 \$2874 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $855 r0 *1 444.495,944.16 sg13_lv_nmos
M$855 VSS \$2874 \$2875 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $859 r0 *1 447.375,944.16 sg13_lv_nmos
M$859 VSS \$2875 \$2876 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $863 r0 *1 450.255,944.16 sg13_lv_nmos
M$863 VSS \$2876 \$2877 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $867 r0 *1 453.135,944.16 sg13_lv_nmos
M$867 VSS \$2877 \$2878 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $871 r0 *1 456.015,944.16 sg13_lv_nmos
M$871 VSS \$2878 \$2879 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $875 r0 *1 461.775,944.16 sg13_lv_nmos
M$875 VSS \$2880 \$2881 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $879 r0 *1 464.595,944.16 sg13_lv_nmos
M$879 VSS \$2881 \$2882 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $887 r0 *1 478.18,943.83 sg13_lv_nmos
M$887 \$2898 \$2942 \$2943 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $888 r0 *1 478.38,942.76 sg13_lv_nmos
M$888 \$2883 \$2882 \$2898 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $889 r0 *1 480.98,942.755 sg13_lv_nmos
M$889 \$2884 \$2882 \$2899 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $890 r0 *1 480.985,943.845 sg13_lv_nmos
M$890 \$2899 \$2943 \$2942 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $891 r0 *1 488.225,943.68 sg13_lv_nmos
M$891 \$2900 \$2932 \$2944 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $892 r0 *1 491.05,943.68 sg13_lv_nmos
M$892 \$2901 \$2944 \$2932 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $893 r0 *1 497.5,943.66 sg13_lv_nmos
M$893 VSS \$2932 \$2933 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $894 r0 *1 498.01,943.61 sg13_lv_nmos
M$894 VSS \$2933 \$2934 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $896 r0 *1 507.67,943.215 sg13_lv_nmos
M$896 \$2892 \$2887 \$2935 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $897 r0 *1 508.18,943.215 sg13_lv_nmos
M$897 \$2935 \$2903 \$2902 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $898 r0 *1 434.915,946.5 sg13_lv_nmos
M$898 VSS \$3013 \$2930 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $900 r0 *1 436.835,946.5 sg13_lv_nmos
M$900 VSS \$2930 \$2981 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $902 r0 *1 438.7,944.185 sg13_lv_nmos
M$902 \$2940 \$2931 \$2873 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $904 r0 *1 439.73,944.185 sg13_lv_nmos
M$904 \$2940 \$2930 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $906 r0 *1 438.7,946.475 sg13_lv_nmos
M$906 \$2982 \$2981 \$2991 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $908 r0 *1 439.73,946.475 sg13_lv_nmos
M$908 \$2982 \$2879 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $910 r0 *1 441.615,946.5 sg13_lv_nmos
M$910 VSS \$2991 \$2983 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $914 r0 *1 444.495,946.5 sg13_lv_nmos
M$914 VSS \$2983 \$2984 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $918 r0 *1 447.375,946.5 sg13_lv_nmos
M$918 VSS \$2984 \$2985 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $922 r0 *1 450.255,946.5 sg13_lv_nmos
M$922 VSS \$2985 \$2986 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $926 r0 *1 453.135,946.5 sg13_lv_nmos
M$926 VSS \$2986 \$2987 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $930 r0 *1 456.015,946.5 sg13_lv_nmos
M$930 VSS \$2987 \$2931 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $934 r0 *1 458.97,946.475 sg13_lv_nmos
M$934 \$2988 \$2931 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $936 r0 *1 460,946.475 sg13_lv_nmos
M$936 \$2988 \$2986 \$2992 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $938 r0 *1 458.97,944.185 sg13_lv_nmos
M$938 \$2941 \$2879 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $940 r0 *1 460,944.185 sg13_lv_nmos
M$940 \$2941 \$2877 \$2880 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $942 r0 *1 461.775,946.5 sg13_lv_nmos
M$942 VSS \$2992 \$2989 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $946 r0 *1 464.595,946.5 sg13_lv_nmos
M$946 VSS \$2989 \$2863 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $954 r0 *1 436.35,962.305 sg13_lv_nmos
M$954 VSS \$2863 \$3053 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $955 r0 *1 437.44,962.4 sg13_lv_nmos
M$955 VSS \$2897 \$3054 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $956 r0 *1 438.29,962.305 sg13_lv_nmos
M$956 VSS \$2882 \$3068 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $957 r0 *1 438.6,962.305 sg13_lv_nmos
M$957 \$3068 \$3054 \$3055 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $958 r0 *1 439.93,962.465 sg13_lv_nmos
M$958 \$3056 \$2882 \$3070 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $959 r0 *1 440.44,962.465 sg13_lv_nmos
M$959 VSS \$2897 \$3070 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $960 r0 *1 440.95,962.415 sg13_lv_nmos
M$960 VSS \$3056 \$3057 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $961 r0 *1 445.76,966.03 sg13_lv_nmos
M$961 PAD|VLO \$3057 \$3093 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $962 r0 *1 448.175,966.09 sg13_lv_nmos
M$962 \$3093 \$2863 CORE$12 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $963 r0 *1 454.2,965.645 sg13_lv_nmos
M$963 VSS \$3099 \$3099 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $964 r0 *1 453.855,962.755 sg13_lv_nmos
M$964 \$3099 \$2987 \$3058 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $965 r0 *1 454.365,962.755 sg13_lv_nmos
M$965 \$3058 \$2882 \$3046 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $966 r0 *1 458.575,965.63 sg13_lv_nmos
M$966 VSS \$3047 \$3048 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $967 r0 *1 458.255,962.735 sg13_lv_nmos
M$967 \$3047 \$2863 \$3046 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $968 r0 *1 458.765,962.735 sg13_lv_nmos
M$968 \$3046 \$173 \$3048 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $969 r0 *1 465.43,962.305 sg13_lv_nmos
M$969 VSS \$2882 \$3059 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $970 r0 *1 466.52,962.4 sg13_lv_nmos
M$970 VSS \$2934 \$3060 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $971 r0 *1 467.37,962.305 sg13_lv_nmos
M$971 VSS \$2863 \$3074 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $972 r0 *1 467.68,962.305 sg13_lv_nmos
M$972 \$3074 \$3060 \$3061 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $973 r0 *1 469.01,962.465 sg13_lv_nmos
M$973 \$3062 \$2863 \$3076 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $974 r0 *1 469.52,962.465 sg13_lv_nmos
M$974 VSS \$2934 \$3076 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $975 r0 *1 470.03,962.415 sg13_lv_nmos
M$975 VSS \$3062 \$3063 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $976 r0 *1 474.84,966.03 sg13_lv_nmos
M$976 PAD|VLO \$3063 \$3094 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $977 r0 *1 477.255,966.09 sg13_lv_nmos
M$977 \$3094 \$2882 \$3048 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $978 r0 *1 483.28,965.645 sg13_lv_nmos
M$978 VSS \$3100 \$3100 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $979 r0 *1 482.935,962.755 sg13_lv_nmos
M$979 \$3100 \$2878 \$3064 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $980 r0 *1 483.445,962.755 sg13_lv_nmos
M$980 \$3064 \$2863 \$3065 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $981 r0 *1 487.655,965.63 sg13_lv_nmos
M$981 VSS \$3049 \$3050 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $982 r0 *1 487.335,962.735 sg13_lv_nmos
M$982 \$3049 \$2882 \$3065 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $983 r0 *1 487.845,962.735 sg13_lv_nmos
M$983 \$3065 \$173 \$3050 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $984 r0 *1 515.91,947.59 sg13_lv_nmos
M$984 VSS \$2897 \$3150 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $986 r0 *1 1060.995,997.48 sg13_lv_nmos
M$986 \$3148 \$3150 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $987 r0 *1 1060.995,1000.99 sg13_lv_nmos
M$987 \$3176 \$3150 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $988 r0 *1 700.255,1060.995 sg13_lv_nmos
M$988 \$1474 \$3240 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $989 r0 *1 800.255,1060.995 sg13_lv_nmos
M$989 \$2651 \$3241 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $990 r0 *1 900.255,1060.995 sg13_lv_nmos
M$990 \$3013 \$3242 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $991 r0 *1 501.765,239.055 sg13_hv_nmos
M$991 VSS CORE \$178 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $992 r0 *1 701.765,239.055 sg13_hv_nmos
M$992 VSS CORE$1 \$179 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $993 r0 *1 801.765,239.055 sg13_hv_nmos
M$993 VSS CORE$2 \$180 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $994 r0 *1 901.765,239.055 sg13_hv_nmos
M$994 VSS CORE$3 \$181 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $995 r0 *1 90.95,285.52 sg13_hv_nmos
M$995 VSS \$219 IN6|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1015 r0 *1 1209.05,294.58 sg13_hv_nmos
M$1015 VSS \$249 OUT6 VSS sg13_hv_nmos W=35.199999999999996 L=0.5999999999999999
* device instance $1023 r0 *1 1064.68,297.64 sg13_hv_nmos
M$1023 \$231 dout VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1024 r0 *1 1064.68,298.47 sg13_hv_nmos
M$1024 VSS \$230 \$241 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1025 r0 *1 1064.68,299.81 sg13_hv_nmos
M$1025 VSS \$241 \$249 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1026 r0 *1 1064.68,301.15 sg13_hv_nmos
M$1026 \$269 dout VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1027 r0 *1 1064.68,301.98 sg13_hv_nmos
M$1027 VSS \$268 \$287 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1028 r0 *1 1064.68,303.32 sg13_hv_nmos
M$1028 VSS \$287 \$209 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1029 r0 *1 90.95,385.52 sg13_hv_nmos
M$1029 VSS \$609 IN5|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1049 r0 *1 1209.05,394.58 sg13_hv_nmos
M$1049 VSS \$672 OUT5 VSS sg13_hv_nmos W=35.199999999999996 L=0.5999999999999999
* device instance $1057 r0 *1 1064.68,397.64 sg13_hv_nmos
M$1057 \$644 \$645 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1058 r0 *1 1064.68,398.47 sg13_hv_nmos
M$1058 VSS \$643 \$665 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1059 r0 *1 1064.68,399.81 sg13_hv_nmos
M$1059 VSS \$665 \$672 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1060 r0 *1 1064.68,401.15 sg13_hv_nmos
M$1060 \$688 \$645 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1061 r0 *1 1064.68,401.98 sg13_hv_nmos
M$1061 VSS \$687 \$698 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1062 r0 *1 1064.68,403.32 sg13_hv_nmos
M$1062 VSS \$698 \$599 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1063 r0 *1 90.95,485.52 sg13_hv_nmos
M$1063 VSS \$1073 IN4|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1083 r0 *1 1209.05,494.58 sg13_hv_nmos
M$1083 VSS \$1100 OUT4 VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999999
* device instance $1091 r0 *1 1064.68,497.64 sg13_hv_nmos
M$1091 \$1084 \$1085 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1092 r0 *1 1064.68,498.47 sg13_hv_nmos
M$1092 VSS \$1083 \$1097 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1093 r0 *1 1064.68,499.81 sg13_hv_nmos
M$1093 VSS \$1097 \$1100 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1094 r0 *1 1064.68,501.15 sg13_hv_nmos
M$1094 \$1112 \$1085 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1095 r0 *1 1064.68,501.98 sg13_hv_nmos
M$1095 VSS \$1111 \$1119 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1096 r0 *1 1064.68,503.32 sg13_hv_nmos
M$1096 VSS \$1119 \$1063 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1097 r0 *1 90.95,585.52 sg13_hv_nmos
M$1097 VSS \$1466 PAD|VLO VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1117 r0 *1 1139.21,663.22 sg13_hv_nmos
M$1117 VSS \$1802 \$1803 VSS sg13_hv_nmos W=108.0 L=0.5
* device instance $1123 r0 *1 1139.21,673 sg13_hv_nmos
M$1123 VSS \$1802 VSS VSS sg13_hv_nmos W=126.0 L=9.5
* device instance $1143 r0 *1 1194.53,668.155 sg13_hv_nmos
M$1143 VSS \$1803 IOVDD VSS sg13_hv_nmos W=756.7999999999977
+ L=0.5999999999999999
* device instance $1315 r0 *1 90.95,685.52 sg13_hv_nmos
M$1315 VSS \$1809 PAD|VHI VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1335 r0 *1 90.95,785.52 sg13_hv_nmos
M$1335 VSS \$1899 IN3|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1355 r0 *1 1209.05,794.58 sg13_hv_nmos
M$1355 VSS \$1926 OUT3 VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999999
* device instance $1363 r0 *1 1064.68,797.64 sg13_hv_nmos
M$1363 \$1910 \$1911 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1364 r0 *1 1064.68,798.47 sg13_hv_nmos
M$1364 VSS \$1909 \$1923 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1365 r0 *1 1064.68,799.81 sg13_hv_nmos
M$1365 VSS \$1923 \$1926 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1366 r0 *1 1064.68,801.15 sg13_hv_nmos
M$1366 \$1938 \$1911 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1367 r0 *1 1064.68,801.98 sg13_hv_nmos
M$1367 VSS \$1937 \$1945 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1368 r0 *1 1064.68,803.32 sg13_hv_nmos
M$1368 VSS \$1945 \$1889 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1369 r0 *1 522.935,859.567 sg13_hv_nmos
M$1369 \$2544 \$2544 VSS VSS sg13_hv_nmos W=33.0 L=0.9
* device instance $1377 r0 *1 542.43,859.567 sg13_hv_nmos
M$1377 \$2546 \$2544 VSS VSS sg13_hv_nmos W=33.0 L=0.9
* device instance $1385 r0 *1 507.575,859.662 sg13_hv_nmos
M$1385 \$2545 \$2544 VSS VSS sg13_hv_nmos W=33.0 L=0.9
* device instance $1393 r0 *1 518.315,858.145 sg13_hv_nmos
M$1393 VSS \$2545 \$2619 VSS sg13_hv_nmos W=1.0 L=0.44999999999999996
* device instance $1394 r0 *1 507.575,870.8 sg13_hv_nmos
M$1394 \$2592 \$2544 \$2619 VSS sg13_hv_nmos W=178.00000000000006
+ L=0.8999999999999999
* device instance $1414 r0 *1 90.95,885.52 sg13_hv_nmos
M$1414 VSS \$2706 IN2|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1434 r0 *1 541.31,863.82 sg13_hv_nmos
M$1434 \$2560 PAD|VLDO \$2546 VSS sg13_hv_nmos W=136.5 L=0.9
* device instance $1448 r0 *1 552.54,863.82 sg13_hv_nmos
M$1448 \$2126 CORE$10 \$2546 VSS sg13_hv_nmos W=136.5 L=0.9
* device instance $1462 r0 *1 1064.68,901.15 sg13_hv_nmos
M$1462 \$2801 \$2391 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1463 r0 *1 1064.68,901.98 sg13_hv_nmos
M$1463 VSS \$2800 \$2808 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1464 r0 *1 1064.68,903.32 sg13_hv_nmos
M$1464 VSS \$2808 \$2683 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1465 r0 *1 1064.68,899.81 sg13_hv_nmos
M$1465 VSS \$2783 \$2789 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1466 r0 *1 1064.68,897.64 sg13_hv_nmos
M$1466 \$2774 \$2391 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1467 r0 *1 1064.68,898.47 sg13_hv_nmos
M$1467 VSS \$2773 \$2783 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1468 r0 *1 1209.05,894.58 sg13_hv_nmos
M$1468 VSS \$2789 OUT2 VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999999
* device instance $1476 r0 *1 90.95,985.52 sg13_hv_nmos
M$1476 VSS \$3138 IN1|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1496 r0 *1 1209.05,994.58 sg13_hv_nmos
M$1496 VSS \$3165 OUT1 VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999999
* device instance $1504 r0 *1 1064.68,997.64 sg13_hv_nmos
M$1504 \$3149 \$3150 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1505 r0 *1 1064.68,998.47 sg13_hv_nmos
M$1505 VSS \$3148 \$3159 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1506 r0 *1 1064.68,999.81 sg13_hv_nmos
M$1506 VSS \$3159 \$3165 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1507 r0 *1 1064.68,1001.15 sg13_hv_nmos
M$1507 \$3177 \$3150 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1508 r0 *1 1064.68,1001.98 sg13_hv_nmos
M$1508 VSS \$3176 \$3184 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1509 r0 *1 1064.68,1003.32 sg13_hv_nmos
M$1509 VSS \$3184 \$3129 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1510 r0 *1 701.765,1060.945 sg13_hv_nmos
M$1510 VSS CORE$13 \$3240 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $1511 r0 *1 801.765,1060.945 sg13_hv_nmos
M$1511 VSS CORE$14 \$3241 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $1512 r0 *1 901.765,1060.945 sg13_hv_nmos
M$1512 VSS CORE$15 \$3242 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $1513 r0 *1 263.22,1139.21 sg13_hv_nmos
M$1513 VSS \$3368 \$3309 VSS sg13_hv_nmos W=108.0 L=0.5
* device instance $1519 r0 *1 273,1139.21 sg13_hv_nmos
M$1519 VSS \$3368 VSS VSS sg13_hv_nmos W=126.0 L=9.5
* device instance $1526 r0 *1 563.22,1139.21 sg13_hv_nmos
M$1526 VSS \$3369 \$3310 VSS sg13_hv_nmos W=108.0 L=0.5
* device instance $1532 r0 *1 573,1139.21 sg13_hv_nmos
M$1532 VSS \$3369 VSS VSS sg13_hv_nmos W=126.0 L=9.5
* device instance $1539 r0 *1 963.22,1139.21 sg13_hv_nmos
M$1539 VSS \$3370 \$3311 VSS sg13_hv_nmos W=108.0 L=0.5
* device instance $1545 r0 *1 973,1139.21 sg13_hv_nmos
M$1545 VSS \$3370 VSS VSS sg13_hv_nmos W=126.0 L=9.5
* device instance $1591 r0 *1 268.155,1194.53 sg13_hv_nmos
M$1591 VSS \$3309 AVDD VSS sg13_hv_nmos W=756.7999999999977 L=0.5999999999999999
* device instance $1634 r0 *1 568.155,1194.53 sg13_hv_nmos
M$1634 VSS \$3310 IOVDD VSS sg13_hv_nmos W=756.7999999999977
+ L=0.5999999999999999
* device instance $1677 r0 *1 968.155,1194.53 sg13_hv_nmos
M$1677 VSS \$3311 VDD VSS sg13_hv_nmos W=756.7999999999977 L=0.5999999999999999
* device instance $2021 r0 *1 385.52,1209.05 sg13_hv_nmos
M$2021 VSS \$3440 PAD|VREF VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $2041 r0 *1 485.52,1209.05 sg13_hv_nmos
M$2041 VSS \$3441 PAD|VLDO VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $2147 r0 *1 500.255,243.995 sg13_lv_pmos
M$2147 \$173 \$178 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2148 r0 *1 700.255,243.995 sg13_lv_pmos
M$2148 \$174 \$179 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2149 r0 *1 800.255,243.995 sg13_lv_pmos
M$2149 \$175 \$180 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2150 r0 *1 900.255,243.995 sg13_lv_pmos
M$2150 \$176 \$181 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2151 r0 *1 1056.005,297.48 sg13_lv_pmos
M$2151 \$230 dout VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2152 r0 *1 431.875,302.8 sg13_lv_pmos
M$2152 VDD \$283 \$270 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2154 r0 *1 432.905,302.8 sg13_lv_pmos
M$2154 VDD \$374 \$270 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2156 r0 *1 434.755,302.8 sg13_lv_pmos
M$2156 VDD \$284 \$263 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2158 r0 *1 435.785,302.8 sg13_lv_pmos
M$2158 VDD \$324 \$263 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2160 r0 *1 437.56,302.8 sg13_lv_pmos
M$2160 VDD \$270 \$264 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2164 r0 *1 440.44,302.8 sg13_lv_pmos
M$2164 VDD \$263 \$265 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2168 r0 *1 443.26,302.8 sg13_lv_pmos
M$2168 VDD \$264 \$266 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2176 r0 *1 448.06,302.8 sg13_lv_pmos
M$2176 VDD \$265 \$267 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2184 r0 *1 1056.005,300.99 sg13_lv_pmos
M$2184 \$268 dout VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2185 r0 *1 431.075,307.485 sg13_lv_pmos
M$2185 VDD \$176 \$319 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2187 r0 *1 433.06,307.485 sg13_lv_pmos
M$2187 VDD \$319 \$331 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2189 r0 *1 434.09,307.485 sg13_lv_pmos
M$2189 VDD \$283 \$331 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2191 r0 *1 435.865,307.485 sg13_lv_pmos
M$2191 VDD \$331 \$321 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2195 r0 *1 438.745,307.485 sg13_lv_pmos
M$2195 VDD \$321 \$322 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2199 r0 *1 441.625,307.485 sg13_lv_pmos
M$2199 VDD \$322 \$323 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2203 r0 *1 444.505,307.485 sg13_lv_pmos
M$2203 VDD \$323 \$324 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2207 r0 *1 447.385,307.485 sg13_lv_pmos
M$2207 VDD \$324 \$325 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2211 r0 *1 450.265,307.485 sg13_lv_pmos
M$2211 VDD \$325 \$284 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2215 r0 *1 456.8,304.885 sg13_lv_pmos
M$2215 VDD \$267 \$291 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2216 r0 *1 457.97,305.01 sg13_lv_pmos
M$2216 VDD \$266 \$294 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2217 r0 *1 458.48,305.01 sg13_lv_pmos
M$2217 VDD \$247 \$294 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2218 r0 *1 458.99,304.87 sg13_lv_pmos
M$2218 VDD \$294 \$295 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2219 r0 *1 460.28,304.73 sg13_lv_pmos
M$2219 \$296 \$247 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2220 r0 *1 460.82,304.87 sg13_lv_pmos
M$2220 VDD \$266 \$292 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2221 r0 *1 461.33,304.87 sg13_lv_pmos
M$2221 \$292 \$296 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2222 r0 *1 431.04,312.135 sg13_lv_pmos
M$2222 VDD \$319 \$368 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2224 r0 *1 433.025,312.135 sg13_lv_pmos
M$2224 VDD \$284 \$370 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2226 r0 *1 434.055,312.135 sg13_lv_pmos
M$2226 VDD \$368 \$370 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2228 r0 *1 435.83,312.135 sg13_lv_pmos
M$2228 VDD \$370 \$371 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2232 r0 *1 438.71,312.135 sg13_lv_pmos
M$2232 VDD \$371 \$372 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2236 r0 *1 441.59,312.135 sg13_lv_pmos
M$2236 VDD \$372 \$373 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2240 r0 *1 444.47,312.135 sg13_lv_pmos
M$2240 VDD \$373 \$374 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2244 r0 *1 447.35,312.135 sg13_lv_pmos
M$2244 VDD \$374 \$375 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2248 r0 *1 450.23,312.135 sg13_lv_pmos
M$2248 VDD \$375 \$283 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2252 r0 *1 457.62,310.765 sg13_lv_pmos
M$2252 \$347 \$292 PAD|VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2253 r0 *1 460.105,309.515 sg13_lv_pmos
M$2253 \$347 \$291 \$346 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2256 r0 *1 431.695,323.31 sg13_lv_pmos
M$2256 VDD \$266 \$442 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2257 r0 *1 432.865,323.435 sg13_lv_pmos
M$2257 VDD \$267 \$446 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2258 r0 *1 433.375,323.435 sg13_lv_pmos
M$2258 VDD \$439 \$446 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2259 r0 *1 433.885,323.295 sg13_lv_pmos
M$2259 VDD \$446 \$443 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2260 r0 *1 435.175,323.155 sg13_lv_pmos
M$2260 \$447 \$439 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2261 r0 *1 435.715,323.295 sg13_lv_pmos
M$2261 VDD \$267 \$444 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2262 r0 *1 436.225,323.295 sg13_lv_pmos
M$2262 \$444 \$447 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2263 r0 *1 451.11,327.385 sg13_lv_pmos
M$2263 VDD \$266 \$467 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2264 r0 *1 452.55,327.385 sg13_lv_pmos
M$2264 VDD \$173 \$493 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2265 r0 *1 454.96,327.385 sg13_lv_pmos
M$2265 VDD \$546 \$494 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2266 r0 *1 453.94,327.37 sg13_lv_pmos
M$2266 VDD \$494 \$247 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2268 r0 *1 461.43,327.36 sg13_lv_pmos
M$2268 \$481 \$463 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2269 r0 *1 462.155,327.36 sg13_lv_pmos
M$2269 VDD \$266 \$463 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2270 r0 *1 465.395,311.56 sg13_lv_pmos
M$2270 AVDD \$297 \$297 AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2274 r0 *1 469.615,311.56 sg13_lv_pmos
M$2274 AVDD \$272 \$271 AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2278 r0 *1 468.43,327.37 sg13_lv_pmos
M$2278 VDD \$473 \$439 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2280 r0 *1 470.55,327.37 sg13_lv_pmos
M$2280 VDD \$439 dout VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2282 r0 *1 435,327.94 sg13_lv_pmos
M$2282 \$480 \$442 CORE$4 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2285 r0 *1 456.085,327.12 sg13_lv_pmos
M$2285 VDD \$546 \$468 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2286 r0 *1 456.595,327.12 sg13_lv_pmos
M$2286 VDD \$493 \$468 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2287 r0 *1 457.045,327.41 sg13_lv_pmos
M$2287 VDD \$495 \$462 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2288 r0 *1 458.095,327.485 sg13_lv_pmos
M$2288 \$495 \$493 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2289 r0 *1 458.83,327.485 sg13_lv_pmos
M$2289 VDD \$462 \$511 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2290 r0 *1 459.22,327.485 sg13_lv_pmos
M$2290 \$511 \$463 \$495 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2291 r0 *1 459.73,327.485 sg13_lv_pmos
M$2291 \$495 \$481 \$468 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2292 r0 *1 464.285,327.105 sg13_lv_pmos
M$2292 \$482 \$481 \$504 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2293 r0 *1 464.665,327.105 sg13_lv_pmos
M$2293 \$504 \$471 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2294 r0 *1 465.275,327.105 sg13_lv_pmos
M$2294 VDD \$493 \$471 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2295 r0 *1 465.785,327.105 sg13_lv_pmos
M$2295 VDD \$482 \$471 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2296 r0 *1 467.345,327.21 sg13_lv_pmos
M$2296 VDD \$482 \$473 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2297 r0 *1 466.325,327.27 sg13_lv_pmos
M$2297 VDD \$482 \$472 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2299 r0 *1 463.59,327.395 sg13_lv_pmos
M$2299 \$462 \$463 \$482 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2300 r0 *1 432.515,329.19 sg13_lv_pmos
M$2300 \$480 \$444 PAD|VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2301 r0 *1 440.29,329.985 sg13_lv_pmos
M$2301 AVDD \$448 \$448 AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2305 r0 *1 444.51,329.985 sg13_lv_pmos
M$2305 AVDD \$440 \$346 AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2309 r0 *1 460.335,334.225 sg13_lv_pmos
M$2309 AVDD \$267 \$543 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2310 r0 *1 460.845,334.225 sg13_lv_pmos
M$2310 \$543 \$544 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2311 r0 *1 463.38,334.225 sg13_lv_pmos
M$2311 AVDD \$543 \$544 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2312 r0 *1 463.89,334.225 sg13_lv_pmos
M$2312 \$544 \$267 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2313 r0 *1 467.145,334.24 sg13_lv_pmos
M$2313 VDD \$544 \$545 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2314 r0 *1 467.655,334.24 sg13_lv_pmos
M$2314 \$545 \$546 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2315 r0 *1 470.18,334.24 sg13_lv_pmos
M$2315 VDD \$545 \$546 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2316 r0 *1 470.69,334.24 sg13_lv_pmos
M$2316 \$546 \$543 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2317 r0 *1 458.31,333.385 sg13_lv_pmos
M$2317 \$526 \$467 \$271 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2320 r0 *1 464.23,395.26 sg13_lv_pmos
M$2320 \$623 \$625 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2321 r0 *1 464.74,395.4 sg13_lv_pmos
M$2321 VDD \$645 \$625 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2322 r0 *1 465.25,395.4 sg13_lv_pmos
M$2322 \$625 \$693 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2323 r0 *1 476.37,395.4 sg13_lv_pmos
M$2323 VDD \$652 \$626 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2324 r0 *1 476.88,395.4 sg13_lv_pmos
M$2324 VDD \$627 \$626 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2325 r0 *1 477.39,395.26 sg13_lv_pmos
M$2325 VDD \$626 \$624 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2326 r0 *1 463.96,399.38 sg13_lv_pmos
M$2326 \$632 \$653 CORE$5 AVDD sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2330 r0 *1 476.13,399.38 sg13_lv_pmos
M$2330 \$659 \$654 \$799 AVDD sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2334 r0 *1 1056.005,397.48 sg13_lv_pmos
M$2334 \$643 \$645 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2335 r0 *1 1056.005,400.99 sg13_lv_pmos
M$2335 \$687 \$645 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2336 r0 *1 466.18,407.01 sg13_lv_pmos
M$2336 PAD|VHI \$711 \$632 AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2337 r0 *1 475.44,407.01 sg13_lv_pmos
M$2337 \$659 \$712 PAD|VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2338 r0 *1 462.07,407.38 sg13_lv_pmos
M$2338 \$721 \$645 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2339 r0 *1 462.61,407.52 sg13_lv_pmos
M$2339 VDD \$693 \$711 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2340 r0 *1 463.12,407.52 sg13_lv_pmos
M$2340 \$711 \$721 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2341 r0 *1 479.55,407.38 sg13_lv_pmos
M$2341 VDD \$627 \$722 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2342 r0 *1 478.5,407.52 sg13_lv_pmos
M$2342 VDD \$722 \$712 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2343 r0 *1 479.01,407.52 sg13_lv_pmos
M$2343 \$712 \$652 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2344 r0 *1 441.985,411.265 sg13_lv_pmos
M$2344 \$696 \$696 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2348 r0 *1 458.735,407.535 sg13_lv_pmos
M$2348 VDD \$652 \$653 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2349 r0 *1 482.89,407.535 sg13_lv_pmos
M$2349 \$654 \$693 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2350 r0 *1 494,411.265 sg13_lv_pmos
M$2350 \$697 \$697 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2354 r0 *1 441.985,420.81 sg13_lv_pmos
M$2354 \$799 \$615 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2358 r0 *1 494,420.81 sg13_lv_pmos
M$2358 \$795 \$618 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2362 r0 *1 452.73,432.655 sg13_lv_pmos
M$2362 VDD \$879 \$847 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2364 r0 *1 453.76,432.655 sg13_lv_pmos
M$2364 VDD \$888 \$847 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2366 r0 *1 455.995,432.655 sg13_lv_pmos
M$2366 VDD \$847 \$839 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2370 r0 *1 459.41,432.655 sg13_lv_pmos
M$2370 VDD \$839 \$840 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2374 r0 *1 462.645,432.655 sg13_lv_pmos
M$2374 VDD \$840 \$841 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2378 r0 *1 466.17,432.655 sg13_lv_pmos
M$2378 VDD \$841 \$842 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2382 r0 *1 470.03,432.655 sg13_lv_pmos
M$2382 VDD \$842 \$843 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2386 r0 *1 474,432.655 sg13_lv_pmos
M$2386 VDD \$843 \$844 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2390 r0 *1 477.92,432.655 sg13_lv_pmos
M$2390 VDD \$844 \$848 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2392 r0 *1 478.95,432.655 sg13_lv_pmos
M$2392 VDD \$842 \$848 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2394 r0 *1 481.6,432.655 sg13_lv_pmos
M$2394 VDD \$848 \$846 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2398 r0 *1 485,432.655 sg13_lv_pmos
M$2398 VDD \$846 \$693 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2406 r0 *1 446.835,440.625 sg13_lv_pmos
M$2406 VDD \$175 \$879 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2408 r0 *1 449.355,440.625 sg13_lv_pmos
M$2408 VDD \$879 \$880 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2410 r0 *1 452.01,440.625 sg13_lv_pmos
M$2410 VDD \$880 \$882 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2412 r0 *1 453.04,440.625 sg13_lv_pmos
M$2412 VDD \$844 \$882 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2414 r0 *1 455.375,440.625 sg13_lv_pmos
M$2414 VDD \$882 \$883 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2418 r0 *1 459.84,440.625 sg13_lv_pmos
M$2418 VDD \$883 \$884 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2422 r0 *1 463.255,440.625 sg13_lv_pmos
M$2422 VDD \$884 \$885 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2426 r0 *1 466.775,440.625 sg13_lv_pmos
M$2426 VDD \$885 \$886 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2430 r0 *1 470.635,440.625 sg13_lv_pmos
M$2430 VDD \$886 \$887 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2434 r0 *1 474.605,440.625 sg13_lv_pmos
M$2434 VDD \$887 \$888 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2438 r0 *1 478.275,440.625 sg13_lv_pmos
M$2438 VDD \$888 \$890 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2440 r0 *1 479.305,440.625 sg13_lv_pmos
M$2440 VDD \$886 \$890 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2442 r0 *1 481.955,440.625 sg13_lv_pmos
M$2442 VDD \$890 \$891 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2446 r0 *1 485.355,440.625 sg13_lv_pmos
M$2446 VDD \$891 \$652 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2454 r0 *1 448.935,453.235 sg13_lv_pmos
M$2454 \$1014 \$988 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2455 r0 *1 448.935,459.035 sg13_lv_pmos
M$2455 \$1044 \$943 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2456 r0 *1 450.345,448.115 sg13_lv_pmos
M$2456 VDD \$1014 \$973 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2457 r0 *1 449.325,448.1 sg13_lv_pmos
M$2457 VDD \$973 \$627 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2459 r0 *1 452.215,447.85 sg13_lv_pmos
M$2459 VDD \$1014 \$953 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2460 r0 *1 452.725,447.85 sg13_lv_pmos
M$2460 VDD \$946 \$953 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2461 r0 *1 453.175,448.14 sg13_lv_pmos
M$2461 VDD \$974 \$948 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2462 r0 *1 452.375,459.035 sg13_lv_pmos
M$2462 VDD \$1014 \$1044 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2463 r0 *1 452.375,453.235 sg13_lv_pmos
M$2463 VDD \$1044 \$1014 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2464 r0 *1 454.225,448.215 sg13_lv_pmos
M$2464 \$974 \$946 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2465 r0 *1 454.96,448.215 sg13_lv_pmos
M$2465 VDD \$948 \$991 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2466 r0 *1 455.35,448.215 sg13_lv_pmos
M$2466 \$991 \$947 \$974 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2467 r0 *1 455.86,448.215 sg13_lv_pmos
M$2467 \$974 \$984 \$953 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2468 r0 *1 457.56,448.09 sg13_lv_pmos
M$2468 \$984 \$947 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2469 r0 *1 458.285,448.09 sg13_lv_pmos
M$2469 VDD \$652 \$947 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2470 r0 *1 460.415,447.835 sg13_lv_pmos
M$2470 \$956 \$984 \$985 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2471 r0 *1 460.795,447.835 sg13_lv_pmos
M$2471 \$985 \$957 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2472 r0 *1 461.405,447.835 sg13_lv_pmos
M$2472 VDD \$946 \$957 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2473 r0 *1 461.915,447.835 sg13_lv_pmos
M$2473 VDD \$956 \$957 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2474 r0 *1 463.475,447.94 sg13_lv_pmos
M$2474 VDD \$956 \$959 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2475 r0 *1 462.455,448 sg13_lv_pmos
M$2475 VDD \$956 \$958 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2477 r0 *1 459.72,448.125 sg13_lv_pmos
M$2477 \$948 \$947 \$956 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2478 r0 *1 464.56,448.1 sg13_lv_pmos
M$2478 VDD \$959 \$645 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2480 r0 *1 467.715,448.115 sg13_lv_pmos
M$2480 VDD \$173 \$946 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2481 r0 *1 469.15,448.115 sg13_lv_pmos
M$2481 VDD \$652 \$960 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2482 r0 *1 470.98,449.055 sg13_lv_pmos
M$2482 \$795 \$960 \$961 AVDD sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2483 r0 *1 481.57,452.025 sg13_lv_pmos
M$2483 AVDD \$943 \$988 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2484 r0 *1 481.57,446.365 sg13_lv_pmos
M$2484 AVDD \$988 \$943 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2485 r0 *1 486.915,446.365 sg13_lv_pmos
M$2485 \$943 \$693 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2486 r0 *1 486.915,452.025 sg13_lv_pmos
M$2486 \$988 \$693 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2487 r0 *1 1056.005,497.48 sg13_lv_pmos
M$2487 \$1083 \$1085 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2488 r0 *1 1056.005,500.99 sg13_lv_pmos
M$2488 \$1111 \$1085 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2489 r0 *1 484.615,506.085 sg13_lv_pmos
M$2489 VDD \$1133 \$1134 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2490 r0 *1 485.125,506.085 sg13_lv_pmos
M$2490 \$1134 \$1145 \$1135 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2491 r0 *1 485.775,506.415 sg13_lv_pmos
M$2491 \$1135 \$1128 \$1169 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2492 r0 *1 486.11,506.415 sg13_lv_pmos
M$2492 \$1169 \$1136 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2493 r0 *1 486.62,506.415 sg13_lv_pmos
M$2493 VDD \$1122 \$1136 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2494 r0 *1 487.13,506.415 sg13_lv_pmos
M$2494 VDD \$1135 \$1136 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2495 r0 *1 487.69,506.25 sg13_lv_pmos
M$2495 VDD \$1135 \$1137 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2496 r0 *1 489.165,506.39 sg13_lv_pmos
M$2496 VDD \$1135 \$1138 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2497 r0 *1 489.675,506.25 sg13_lv_pmos
M$2497 VDD \$1138 \$1139 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2498 r0 *1 491.89,506.25 sg13_lv_pmos
M$2498 VDD \$1139 \$1085 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2500 r0 *1 497.63,506.265 sg13_lv_pmos
M$2500 VDD \$1204 \$1152 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2501 r0 *1 496.61,506.25 sg13_lv_pmos
M$2501 VDD \$1152 \$1140 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2503 r0 *1 476.78,506.265 sg13_lv_pmos
M$2503 VDD \$1305 \$1131 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2504 r0 *1 480.305,506.31 sg13_lv_pmos
M$2504 \$1145 \$1305 VDD VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2505 r0 *1 480.815,506.31 sg13_lv_pmos
M$2505 VDD \$1145 \$1128 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2506 r0 *1 481.975,506.375 sg13_lv_pmos
M$2506 \$1132 \$1128 \$1133 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2507 r0 *1 482.485,506.375 sg13_lv_pmos
M$2507 \$1133 \$1145 \$1167 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2508 r0 *1 482.86,506.375 sg13_lv_pmos
M$2508 \$1167 \$1134 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2509 r0 *1 483.435,506.375 sg13_lv_pmos
M$2509 VDD \$1122 \$1133 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2510 r0 *1 494.705,506.265 sg13_lv_pmos
M$2510 VDD \$173 \$1122 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2511 r0 *1 478.775,506.6 sg13_lv_pmos
M$2511 VDD \$1204 \$1132 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2512 r0 *1 479.285,506.6 sg13_lv_pmos
M$2512 \$1132 \$1122 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2513 r0 *1 481.4,518.61 sg13_lv_pmos
M$2513 \$1199 \$1243 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2514 r0 *1 482.8,518.61 sg13_lv_pmos
M$2514 AVDD \$1200 \$1199 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2515 r0 *1 484.2,518.61 sg13_lv_pmos
M$2515 \$1200 \$1199 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2516 r0 *1 485.6,518.61 sg13_lv_pmos
M$2516 AVDD \$1243 \$1200 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2517 r0 *1 489.12,508.99 sg13_lv_pmos
M$2517 \$1182 \$1131 \$1183 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2520 r0 *1 488.26,518.61 sg13_lv_pmos
M$2520 \$1203 \$1200 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2521 r0 *1 489.66,518.61 sg13_lv_pmos
M$2521 VDD \$1204 \$1203 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2522 r0 *1 491.06,518.61 sg13_lv_pmos
M$2522 \$1204 \$1203 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2523 r0 *1 492.46,518.61 sg13_lv_pmos
M$2523 VDD \$1199 \$1204 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2524 r0 *1 435.35,517.185 sg13_lv_pmos
M$2524 VDD \$1302 \$1234 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2526 r0 *1 436.38,517.185 sg13_lv_pmos
M$2526 VDD \$1249 \$1234 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2528 r0 *1 438.155,517.185 sg13_lv_pmos
M$2528 VDD \$1234 \$1235 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2532 r0 *1 441.035,517.185 sg13_lv_pmos
M$2532 VDD \$1235 \$1236 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2536 r0 *1 443.915,517.185 sg13_lv_pmos
M$2536 VDD \$1236 \$1237 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2540 r0 *1 446.795,517.185 sg13_lv_pmos
M$2540 VDD \$1237 \$1238 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2544 r0 *1 449.675,517.185 sg13_lv_pmos
M$2544 VDD \$1238 \$1239 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2548 r0 *1 452.555,517.185 sg13_lv_pmos
M$2548 VDD \$1239 \$1240 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2552 r0 *1 455.51,517.185 sg13_lv_pmos
M$2552 VDD \$1240 \$1241 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2554 r0 *1 456.54,517.185 sg13_lv_pmos
M$2554 VDD \$1238 \$1241 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2556 r0 *1 458.315,517.185 sg13_lv_pmos
M$2556 VDD \$1241 \$1242 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2560 r0 *1 461.135,517.185 sg13_lv_pmos
M$2560 VDD \$1242 \$1243 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2568 r0 *1 431.445,522.94 sg13_lv_pmos
M$2568 VDD \$174 \$1249 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2570 r0 *1 432.935,536.78 sg13_lv_pmos
M$2570 \$1352 \$1139 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2571 r0 *1 433.475,536.92 sg13_lv_pmos
M$2571 VDD \$1243 \$1353 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2572 r0 *1 433.985,536.92 sg13_lv_pmos
M$2572 \$1353 \$1352 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2573 r0 *1 433.365,522.94 sg13_lv_pmos
M$2573 VDD \$1249 \$1295 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2575 r0 *1 435.35,522.94 sg13_lv_pmos
M$2575 VDD \$1240 \$1308 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2577 r0 *1 436.38,522.94 sg13_lv_pmos
M$2577 VDD \$1295 \$1308 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2579 r0 *1 438.155,522.94 sg13_lv_pmos
M$2579 VDD \$1308 \$1297 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2583 r0 *1 441.035,522.94 sg13_lv_pmos
M$2583 VDD \$1297 \$1298 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2587 r0 *1 443.915,522.94 sg13_lv_pmos
M$2587 VDD \$1298 \$1299 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2591 r0 *1 446.795,522.94 sg13_lv_pmos
M$2591 VDD \$1299 \$1300 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2595 r0 *1 449.675,522.94 sg13_lv_pmos
M$2595 VDD \$1300 \$1301 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2599 r0 *1 452.555,522.94 sg13_lv_pmos
M$2599 VDD \$1301 \$1302 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2603 r0 *1 455.51,522.94 sg13_lv_pmos
M$2603 VDD \$1302 \$1309 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2605 r0 *1 456.54,522.94 sg13_lv_pmos
M$2605 VDD \$1300 \$1309 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2607 r0 *1 458.315,522.94 sg13_lv_pmos
M$2607 VDD \$1309 \$1304 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2611 r0 *1 461.135,522.94 sg13_lv_pmos
M$2611 VDD \$1304 \$1305 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2619 r0 *1 467.935,536.78 sg13_lv_pmos
M$2619 \$1358 \$1140 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2620 r0 *1 468.475,536.92 sg13_lv_pmos
M$2620 VDD \$1305 \$1359 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2621 r0 *1 468.985,536.92 sg13_lv_pmos
M$2621 \$1359 \$1358 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2622 r0 *1 431.51,536.935 sg13_lv_pmos
M$2622 VDD \$1305 \$1351 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2623 r0 *1 435.785,537.06 sg13_lv_pmos
M$2623 VDD \$1243 \$1354 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2624 r0 *1 436.295,537.06 sg13_lv_pmos
M$2624 VDD \$1139 \$1354 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2625 r0 *1 436.805,536.92 sg13_lv_pmos
M$2625 VDD \$1354 \$1355 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2626 r0 *1 452.575,539.207 sg13_lv_pmos
M$2626 \$1372 \$1377 AVDD AVDD sg13_lv_pmos W=10.5 L=1.5
* device instance $2630 r0 *1 466.51,536.935 sg13_lv_pmos
M$2630 VDD \$1243 \$1357 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2631 r0 *1 470.785,537.06 sg13_lv_pmos
M$2631 VDD \$1305 \$1360 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2632 r0 *1 471.295,537.06 sg13_lv_pmos
M$2632 VDD \$1140 \$1360 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2633 r0 *1 471.805,536.92 sg13_lv_pmos
M$2633 VDD \$1360 \$1361 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2634 r0 *1 487.575,539.207 sg13_lv_pmos
M$2634 \$1182 \$1378 AVDD AVDD sg13_lv_pmos W=10.5 L=1.5
* device instance $2638 r0 *1 440.925,539.222 sg13_lv_pmos
M$2638 \$1356 \$1356 AVDD AVDD sg13_lv_pmos W=10.5 L=1.5
* device instance $2642 r0 *1 475.925,539.222 sg13_lv_pmos
M$2642 \$1189 \$1189 AVDD AVDD sg13_lv_pmos W=10.5 L=1.5
* device instance $2646 r0 *1 434.41,549.415 sg13_lv_pmos
M$2646 \$1401 \$1353 PAD|VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2647 r0 *1 436.765,548.915 sg13_lv_pmos
M$2647 \$1401 \$1351 CORE$6 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2650 r0 *1 469.41,549.415 sg13_lv_pmos
M$2650 \$1402 \$1359 PAD|VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2651 r0 *1 471.765,548.915 sg13_lv_pmos
M$2651 \$1402 \$1357 \$1372 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2654 r0 *1 449.83,598.84 sg13_lv_pmos
M$2654 VDD \$1532 \$1489 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2656 r0 *1 450.86,598.84 sg13_lv_pmos
M$2656 VDD \$1488 \$1489 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2658 r0 *1 452.635,598.84 sg13_lv_pmos
M$2658 VDD \$1489 \$1479 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2662 r0 *1 455.515,598.84 sg13_lv_pmos
M$2662 VDD \$1479 \$1480 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2666 r0 *1 458.395,598.84 sg13_lv_pmos
M$2666 VDD \$1480 \$1481 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2670 r0 *1 461.275,598.84 sg13_lv_pmos
M$2670 VDD \$1481 \$1482 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2674 r0 *1 464.155,598.84 sg13_lv_pmos
M$2674 VDD \$1482 \$1483 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2678 r0 *1 467.035,598.84 sg13_lv_pmos
M$2678 VDD \$1483 \$1484 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2682 r0 *1 469.99,598.84 sg13_lv_pmos
M$2682 VDD \$1484 \$1490 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2684 r0 *1 471.02,598.84 sg13_lv_pmos
M$2684 VDD \$1482 \$1490 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2686 r0 *1 472.795,598.84 sg13_lv_pmos
M$2686 VDD \$1490 \$1486 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2690 r0 *1 475.615,598.84 sg13_lv_pmos
M$2690 VDD \$1486 \$1487 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2698 r0 *1 445.925,604.64 sg13_lv_pmos
M$2698 VDD \$1474 \$1488 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2700 r0 *1 447.845,604.64 sg13_lv_pmos
M$2700 VDD \$1488 \$1524 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2702 r0 *1 449.83,604.64 sg13_lv_pmos
M$2702 VDD \$1484 \$1526 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2704 r0 *1 450.86,604.64 sg13_lv_pmos
M$2704 VDD \$1524 \$1526 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2706 r0 *1 452.635,604.64 sg13_lv_pmos
M$2706 VDD \$1526 \$1527 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2710 r0 *1 455.515,604.64 sg13_lv_pmos
M$2710 VDD \$1527 \$1528 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2714 r0 *1 458.395,604.64 sg13_lv_pmos
M$2714 VDD \$1528 \$1529 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2718 r0 *1 461.275,604.64 sg13_lv_pmos
M$2718 VDD \$1529 \$1530 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2722 r0 *1 464.155,604.64 sg13_lv_pmos
M$2722 VDD \$1530 \$1531 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2726 r0 *1 467.035,604.64 sg13_lv_pmos
M$2726 VDD \$1531 \$1532 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2730 r0 *1 469.99,604.64 sg13_lv_pmos
M$2730 VDD \$1532 \$1534 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2732 r0 *1 471.02,604.64 sg13_lv_pmos
M$2732 VDD \$1530 \$1534 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2734 r0 *1 472.795,604.64 sg13_lv_pmos
M$2734 VDD \$1534 \$1535 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2738 r0 *1 475.615,604.64 sg13_lv_pmos
M$2738 VDD \$1535 \$1536 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2746 r0 *1 433.28,618.09 sg13_lv_pmos
M$2746 VDD \$1536 \$1594 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2747 r0 *1 434.36,617.935 sg13_lv_pmos
M$2747 \$1598 \$1567 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2748 r0 *1 434.9,618.075 sg13_lv_pmos
M$2748 VDD \$1487 \$1595 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2749 r0 *1 435.41,618.075 sg13_lv_pmos
M$2749 \$1595 \$1598 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2750 r0 *1 434.995,621.675 sg13_lv_pmos
M$2750 CORE$9 \$1594 \$1653 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2753 r0 *1 436.85,618.215 sg13_lv_pmos
M$2753 VDD \$1487 \$1603 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2754 r0 *1 437.36,618.215 sg13_lv_pmos
M$2754 VDD \$1567 \$1603 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2755 r0 *1 437.87,618.075 sg13_lv_pmos
M$2755 VDD \$1603 \$1587 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2756 r0 *1 439.97,617.765 sg13_lv_pmos
M$2756 PAD|VHI \$1595 \$1653 AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2757 r0 *1 469.335,618.09 sg13_lv_pmos
M$2757 VDD \$1487 \$1596 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2758 r0 *1 470.415,617.935 sg13_lv_pmos
M$2758 \$1599 \$1568 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2759 r0 *1 470.955,618.075 sg13_lv_pmos
M$2759 VDD \$1536 \$1597 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2760 r0 *1 471.465,618.075 sg13_lv_pmos
M$2760 \$1597 \$1599 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2761 r0 *1 471.05,621.675 sg13_lv_pmos
M$2761 \$1633 \$1596 \$1654 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2764 r0 *1 472.905,618.215 sg13_lv_pmos
M$2764 VDD \$1536 \$1604 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2765 r0 *1 473.415,618.215 sg13_lv_pmos
M$2765 VDD \$1568 \$1604 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2766 r0 *1 473.925,618.075 sg13_lv_pmos
M$2766 VDD \$1604 \$1589 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2767 r0 *1 476.025,617.765 sg13_lv_pmos
M$2767 PAD|VHI \$1597 \$1654 AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2768 r0 *1 505.435,618.205 sg13_lv_pmos
M$2768 VDD \$1536 \$1600 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2769 r0 *1 520.805,621.42 sg13_lv_pmos
M$2769 VDD \$1664 \$1665 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2770 r0 *1 521.315,621.42 sg13_lv_pmos
M$2770 VDD \$1649 \$1665 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2771 r0 *1 521.765,621.71 sg13_lv_pmos
M$2771 VDD \$1680 \$1655 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2772 r0 *1 526.15,621.66 sg13_lv_pmos
M$2772 \$1691 \$1656 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2773 r0 *1 526.875,621.66 sg13_lv_pmos
M$2773 VDD \$1536 \$1656 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2774 r0 *1 529.005,621.405 sg13_lv_pmos
M$2774 \$1666 \$1691 \$1701 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2775 r0 *1 529.385,621.405 sg13_lv_pmos
M$2775 \$1701 \$1658 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2776 r0 *1 529.995,621.405 sg13_lv_pmos
M$2776 VDD \$1649 \$1658 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2777 r0 *1 530.505,621.405 sg13_lv_pmos
M$2777 VDD \$1666 \$1658 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2778 r0 *1 532.065,621.51 sg13_lv_pmos
M$2778 VDD \$1666 \$1660 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2779 r0 *1 531.045,621.57 sg13_lv_pmos
M$2779 VDD \$1666 \$1659 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2781 r0 *1 528.31,621.695 sg13_lv_pmos
M$2781 \$1655 \$1656 \$1666 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2782 r0 *1 533.15,621.67 sg13_lv_pmos
M$2782 VDD \$1660 \$1567 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2784 r0 *1 535.2,621.67 sg13_lv_pmos
M$2784 VDD \$1567 \$1911 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2786 r0 *1 536.99,621.685 sg13_lv_pmos
M$2786 \$1649 \$173 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2787 r0 *1 456.64,625.975 sg13_lv_pmos
M$2787 \$1633 \$1723 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2791 r0 *1 462.64,625.975 sg13_lv_pmos
M$2791 \$1588 \$1588 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2795 r0 *1 492.695,625.975 sg13_lv_pmos
M$2795 \$1634 \$1724 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2799 r0 *1 498.695,625.975 sg13_lv_pmos
M$2799 \$1590 \$1590 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2803 r0 *1 505.15,621.115 sg13_lv_pmos
M$2803 \$1679 \$1600 \$1634 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2806 r0 *1 521.51,632.615 sg13_lv_pmos
M$2806 VDD \$1752 \$1747 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2807 r0 *1 522.815,621.785 sg13_lv_pmos
M$2807 \$1680 \$1649 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2808 r0 *1 523.55,621.785 sg13_lv_pmos
M$2808 VDD \$1655 \$1702 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2809 r0 *1 523.94,621.785 sg13_lv_pmos
M$2809 \$1702 \$1656 \$1680 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2810 r0 *1 524.45,621.785 sg13_lv_pmos
M$2810 \$1680 \$1691 \$1665 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2811 r0 *1 524.18,632.615 sg13_lv_pmos
M$2811 \$1747 \$1664 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2812 r0 *1 528.19,632.615 sg13_lv_pmos
M$2812 VDD \$1747 \$1664 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2813 r0 *1 530.86,632.615 sg13_lv_pmos
M$2813 \$1664 \$1751 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2814 r0 *1 534.455,625.47 sg13_lv_pmos
M$2814 VDD \$1721 \$1568 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2816 r0 *1 534.47,626.49 sg13_lv_pmos
M$2816 VDD \$1664 \$1721 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2817 r0 *1 508.41,633.315 sg13_lv_pmos
M$2817 AVDD \$1487 \$1751 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2818 r0 *1 511.055,633.315 sg13_lv_pmos
M$2818 \$1751 \$1752 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2819 r0 *1 513.41,633.315 sg13_lv_pmos
M$2819 AVDD \$1751 \$1752 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2820 r0 *1 516.045,633.315 sg13_lv_pmos
M$2820 \$1752 \$1487 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2821 r0 *1 1056.005,797.48 sg13_lv_pmos
M$2821 \$1909 \$1911 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2822 r0 *1 1056.005,800.99 sg13_lv_pmos
M$2822 \$1937 \$1911 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2823 r0 *1 633.21,840.21 sg13_lv_pmos
M$2823 PAD|VLDO \$2141 \$2141 PAD|VLDO sg13_lv_pmos W=10.0 L=1.5
* device instance $2825 r0 *1 630.06,845.38 sg13_lv_pmos
M$2825 \$2209 \$2263 \$2174 PAD|VLDO sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2827 r0 *1 622.075,848.775 sg13_lv_pmos
M$2827 PAD|VLDO \$2339 \$2248 PAD|VLDO sg13_lv_pmos W=4.0 L=0.13
* device instance $2829 r0 *1 624.015,848.775 sg13_lv_pmos
M$2829 PAD|VLDO \$2247 \$2248 PAD|VLDO sg13_lv_pmos W=4.0 L=0.13
* device instance $2831 r0 *1 625.955,848.775 sg13_lv_pmos
M$2831 PAD|VLDO \$2248 \$2247 PAD|VLDO sg13_lv_pmos W=4.0 L=0.13
* device instance $2833 r0 *1 627.895,848.775 sg13_lv_pmos
M$2833 PAD|VLDO \$2339 \$2247 PAD|VLDO sg13_lv_pmos W=4.0 L=0.13
* device instance $2835 r0 *1 631.3,848.775 sg13_lv_pmos
M$2835 VDD \$2247 \$2258 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2837 r0 *1 633.24,848.775 sg13_lv_pmos
M$2837 VDD \$2249 \$2258 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2839 r0 *1 635.18,848.775 sg13_lv_pmos
M$2839 VDD \$2258 \$2249 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2841 r0 *1 637.12,848.775 sg13_lv_pmos
M$2841 VDD \$2248 \$2249 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2843 r0 *1 585.345,849.525 sg13_lv_pmos
M$2843 \$2256 \$2335 CORE$11 PAD|VLDO sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2845 r0 *1 586.14,853.855 sg13_lv_pmos
M$2845 PAD|VHI \$2456 \$2256 PAD|VLDO sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2846 r0 *1 592.87,850.555 sg13_lv_pmos
M$2846 PAD|VLDO \$2180 \$2164 PAD|VLDO sg13_lv_pmos W=10.0 L=1.5
* device instance $2848 r0 *1 606.935,849.525 sg13_lv_pmos
M$2848 \$2257 \$2336 \$2164 PAD|VLDO sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2850 r0 *1 607.73,853.855 sg13_lv_pmos
M$2850 PAD|VHI \$2457 \$2257 PAD|VLDO sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2851 r0 *1 614.46,850.555 sg13_lv_pmos
M$2851 PAD|VLDO \$2181 \$2209 PAD|VLDO sg13_lv_pmos W=10.0 L=1.5
* device instance $2853 r0 *1 628.87,853.995 sg13_lv_pmos
M$2853 \$2397 \$2341 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2854 r0 *1 629.595,853.995 sg13_lv_pmos
M$2854 VDD \$2281 \$2341 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2855 r0 *1 620.95,854.02 sg13_lv_pmos
M$2855 VDD \$2281 \$2263 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2856 r0 *1 622.39,854.02 sg13_lv_pmos
M$2856 VDD \$173 \$2385 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2857 r0 *1 635.87,854.005 sg13_lv_pmos
M$2857 VDD \$2390 \$2561 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2859 r0 *1 637.86,854.02 sg13_lv_pmos
M$2859 VDD \$2249 \$2399 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2860 r0 *1 638.37,854.005 sg13_lv_pmos
M$2860 VDD \$2399 \$2562 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2862 r0 *1 640.39,854.005 sg13_lv_pmos
M$2862 VDD \$2561 \$2391 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2864 r0 *1 617.465,865.11 sg13_lv_pmos
M$2864 VDD \$2597 \$2578 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2866 r0 *1 618.495,865.11 sg13_lv_pmos
M$2866 VDD \$2598 \$2578 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2868 r0 *1 620.495,865.11 sg13_lv_pmos
M$2868 VDD \$2578 \$2564 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2872 r0 *1 623.375,865.11 sg13_lv_pmos
M$2872 VDD \$2564 \$2565 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2876 r0 *1 623.525,853.755 sg13_lv_pmos
M$2876 VDD \$2249 \$2386 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2877 r0 *1 624.035,853.755 sg13_lv_pmos
M$2877 VDD \$2385 \$2386 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2878 r0 *1 624.485,854.045 sg13_lv_pmos
M$2878 VDD \$2458 \$2340 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2879 r0 *1 625.535,854.12 sg13_lv_pmos
M$2879 \$2458 \$2385 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2880 r0 *1 626.27,854.12 sg13_lv_pmos
M$2880 VDD \$2340 \$2483 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2881 r0 *1 626.66,854.12 sg13_lv_pmos
M$2881 \$2483 \$2341 \$2458 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2882 r0 *1 627.17,854.12 sg13_lv_pmos
M$2882 \$2458 \$2397 \$2386 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2883 r0 *1 626.255,865.11 sg13_lv_pmos
M$2883 VDD \$2565 \$2566 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2887 r0 *1 629.135,865.11 sg13_lv_pmos
M$2887 VDD \$2566 \$2567 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2891 r0 *1 631.725,853.74 sg13_lv_pmos
M$2891 \$2398 \$2397 \$2474 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2892 r0 *1 632.105,853.74 sg13_lv_pmos
M$2892 \$2474 \$2388 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2893 r0 *1 632.715,853.74 sg13_lv_pmos
M$2893 VDD \$2385 \$2388 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2894 r0 *1 633.225,853.74 sg13_lv_pmos
M$2894 VDD \$2398 \$2388 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2895 r0 *1 634.785,853.845 sg13_lv_pmos
M$2895 VDD \$2398 \$2390 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2896 r0 *1 633.765,853.905 sg13_lv_pmos
M$2896 VDD \$2398 \$2389 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2898 r0 *1 631.03,854.03 sg13_lv_pmos
M$2898 \$2340 \$2341 \$2398 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2899 r0 *1 632.715,865.11 sg13_lv_pmos
M$2899 VDD \$2567 \$2314 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2903 r0 *1 636.295,865.11 sg13_lv_pmos
M$2903 VDD \$2314 \$2568 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2907 r0 *1 640.7,865.11 sg13_lv_pmos
M$2907 VDD \$2568 \$2579 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2909 r0 *1 641.73,865.11 sg13_lv_pmos
M$2909 VDD \$2567 \$2579 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2911 r0 *1 643.75,865.11 sg13_lv_pmos
M$2911 VDD \$2579 \$2570 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2915 r0 *1 646.57,865.11 sg13_lv_pmos
M$2915 VDD \$2570 \$2339 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2923 r0 *1 577.495,865.995 sg13_lv_pmos
M$2923 VDD \$2339 \$2593 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2924 r0 *1 578.005,865.995 sg13_lv_pmos
M$2924 VDD \$2561 \$2593 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2925 r0 *1 578.515,865.855 sg13_lv_pmos
M$2925 VDD \$2593 \$2394 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2926 r0 *1 579.805,865.715 sg13_lv_pmos
M$2926 \$2594 \$2561 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2927 r0 *1 580.345,865.855 sg13_lv_pmos
M$2927 VDD \$2339 \$2456 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2928 r0 *1 580.855,865.855 sg13_lv_pmos
M$2928 \$2456 \$2594 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2929 r0 *1 582.565,865.87 sg13_lv_pmos
M$2929 VDD \$2281 \$2335 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2930 r0 *1 599.085,865.995 sg13_lv_pmos
M$2930 VDD \$2281 \$2595 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2931 r0 *1 599.595,865.995 sg13_lv_pmos
M$2931 VDD \$2562 \$2595 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2932 r0 *1 600.105,865.855 sg13_lv_pmos
M$2932 VDD \$2595 \$2395 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2933 r0 *1 601.395,865.715 sg13_lv_pmos
M$2933 \$2596 \$2562 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2934 r0 *1 601.935,865.855 sg13_lv_pmos
M$2934 VDD \$2281 \$2457 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2935 r0 *1 602.445,865.855 sg13_lv_pmos
M$2935 \$2457 \$2596 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2936 r0 *1 604.155,865.87 sg13_lv_pmos
M$2936 VDD \$2339 \$2336 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2937 r0 *1 613.56,870.785 sg13_lv_pmos
M$2937 VDD \$2651 \$2598 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2939 r0 *1 615.48,870.785 sg13_lv_pmos
M$2939 VDD \$2598 \$2640 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2941 r0 *1 617.465,870.785 sg13_lv_pmos
M$2941 VDD \$2568 \$2642 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2943 r0 *1 618.495,870.785 sg13_lv_pmos
M$2943 VDD \$2640 \$2642 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2945 r0 *1 620.495,870.785 sg13_lv_pmos
M$2945 VDD \$2642 \$2643 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2949 r0 *1 623.375,870.785 sg13_lv_pmos
M$2949 VDD \$2643 \$2644 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2953 r0 *1 626.255,870.785 sg13_lv_pmos
M$2953 VDD \$2644 \$2645 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2957 r0 *1 629.135,870.785 sg13_lv_pmos
M$2957 VDD \$2645 \$2646 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2961 r0 *1 632.715,870.785 sg13_lv_pmos
M$2961 VDD \$2646 \$2647 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2965 r0 *1 636.295,870.785 sg13_lv_pmos
M$2965 VDD \$2647 \$2597 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2969 r0 *1 640.44,870.785 sg13_lv_pmos
M$2969 VDD \$2597 \$2649 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2971 r0 *1 641.47,870.785 sg13_lv_pmos
M$2971 VDD \$2646 \$2649 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2973 r0 *1 643.505,870.785 sg13_lv_pmos
M$2973 VDD \$2649 \$2650 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2977 r0 *1 646.325,870.785 sg13_lv_pmos
M$2977 VDD \$2650 \$2281 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2985 r0 *1 1056.005,897.48 sg13_lv_pmos
M$2985 \$2773 \$2391 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2986 r0 *1 1056.005,900.99 sg13_lv_pmos
M$2986 \$2800 \$2391 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2987 r0 *1 478.37,933.46 sg13_lv_pmos
M$2987 \$2861 \$2859 \$3050 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2990 r0 *1 483.435,934.515 sg13_lv_pmos
M$2990 VDD \$2863 \$2859 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2991 r0 *1 438.7,942.5 sg13_lv_pmos
M$2991 VDD \$2931 \$2873 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2993 r0 *1 439.73,942.5 sg13_lv_pmos
M$2993 VDD \$2930 \$2873 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2995 r0 *1 441.615,942.5 sg13_lv_pmos
M$2995 VDD \$2873 \$2874 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2999 r0 *1 444.495,942.5 sg13_lv_pmos
M$2999 VDD \$2874 \$2875 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3003 r0 *1 447.375,942.5 sg13_lv_pmos
M$3003 VDD \$2875 \$2876 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3007 r0 *1 450.255,942.5 sg13_lv_pmos
M$3007 VDD \$2876 \$2877 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3011 r0 *1 453.135,942.5 sg13_lv_pmos
M$3011 VDD \$2877 \$2878 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3015 r0 *1 456.015,942.5 sg13_lv_pmos
M$3015 VDD \$2878 \$2879 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3019 r0 *1 458.97,942.5 sg13_lv_pmos
M$3019 VDD \$2879 \$2880 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3021 r0 *1 460,942.5 sg13_lv_pmos
M$3021 VDD \$2877 \$2880 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3023 r0 *1 461.775,942.5 sg13_lv_pmos
M$3023 VDD \$2880 \$2881 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3027 r0 *1 464.595,942.5 sg13_lv_pmos
M$3027 VDD \$2881 \$2882 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $3035 r0 *1 434.905,948.16 sg13_lv_pmos
M$3035 VDD \$3013 \$2930 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3037 r0 *1 436.825,948.16 sg13_lv_pmos
M$3037 VDD \$2930 \$2981 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3039 r0 *1 438.7,948.16 sg13_lv_pmos
M$3039 VDD \$2981 \$2991 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3041 r0 *1 439.73,948.16 sg13_lv_pmos
M$3041 VDD \$2879 \$2991 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3043 r0 *1 441.615,948.16 sg13_lv_pmos
M$3043 VDD \$2991 \$2983 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3047 r0 *1 444.495,948.16 sg13_lv_pmos
M$3047 VDD \$2983 \$2984 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3051 r0 *1 447.375,948.16 sg13_lv_pmos
M$3051 VDD \$2984 \$2985 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3055 r0 *1 450.255,948.16 sg13_lv_pmos
M$3055 VDD \$2985 \$2986 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3059 r0 *1 453.135,948.16 sg13_lv_pmos
M$3059 VDD \$2986 \$2987 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3063 r0 *1 456.015,948.16 sg13_lv_pmos
M$3063 VDD \$2987 \$2931 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3067 r0 *1 458.97,948.16 sg13_lv_pmos
M$3067 VDD \$2931 \$2992 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3069 r0 *1 460,948.16 sg13_lv_pmos
M$3069 VDD \$2986 \$2992 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3071 r0 *1 461.775,948.16 sg13_lv_pmos
M$3071 VDD \$2992 \$2989 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3075 r0 *1 464.595,948.16 sg13_lv_pmos
M$3075 VDD \$2989 \$2863 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $3083 r0 *1 477.19,946.75 sg13_lv_pmos
M$3083 \$2943 \$2882 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3084 r0 *1 477.19,945.32 sg13_lv_pmos
M$3084 \$2943 \$2942 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3085 r0 *1 481.99,945.32 sg13_lv_pmos
M$3085 \$2942 \$2882 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3086 r0 *1 481.99,946.75 sg13_lv_pmos
M$3086 \$2942 \$2943 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3087 r0 *1 487.085,945.32 sg13_lv_pmos
M$3087 \$2944 \$2932 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3088 r0 *1 487.085,946.75 sg13_lv_pmos
M$3088 \$2944 \$2942 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3089 r0 *1 492.11,946.735 sg13_lv_pmos
M$3089 \$2932 \$2944 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3090 r0 *1 492.11,945.305 sg13_lv_pmos
M$3090 \$2932 \$2943 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3091 r0 *1 497.5,945.285 sg13_lv_pmos
M$3091 VDD \$2932 \$2933 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $3092 r0 *1 498.01,945.27 sg13_lv_pmos
M$3092 VDD \$2933 \$2934 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3094 r0 *1 503.36,944.28 sg13_lv_pmos
M$3094 VDD \$173 \$2885 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3095 r0 *1 504.495,944.015 sg13_lv_pmos
M$3095 VDD \$2932 \$2892 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3096 r0 *1 505.005,944.015 sg13_lv_pmos
M$3096 VDD \$2885 \$2892 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3097 r0 *1 505.455,944.305 sg13_lv_pmos
M$3097 VDD \$2935 \$2886 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $3098 r0 *1 506.505,944.38 sg13_lv_pmos
M$3098 \$2935 \$2885 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3099 r0 *1 507.24,944.38 sg13_lv_pmos
M$3099 VDD \$2886 \$2962 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3100 r0 *1 507.63,944.38 sg13_lv_pmos
M$3100 \$2962 \$2887 \$2935 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3101 r0 *1 508.14,944.38 sg13_lv_pmos
M$3101 \$2935 \$2903 \$2892 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3102 r0 *1 509.84,944.255 sg13_lv_pmos
M$3102 \$2903 \$2887 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3103 r0 *1 510.565,944.255 sg13_lv_pmos
M$3103 VDD \$2863 \$2887 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3104 r0 *1 512.695,944 sg13_lv_pmos
M$3104 \$2904 \$2903 \$2951 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3105 r0 *1 513.075,944 sg13_lv_pmos
M$3105 \$2951 \$2894 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3106 r0 *1 513.685,944 sg13_lv_pmos
M$3106 VDD \$2885 \$2894 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3107 r0 *1 514.195,944 sg13_lv_pmos
M$3107 VDD \$2904 \$2894 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3108 r0 *1 515.755,944.105 sg13_lv_pmos
M$3108 VDD \$2904 \$2896 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $3109 r0 *1 514.735,944.165 sg13_lv_pmos
M$3109 VDD \$2904 \$2895 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3111 r0 *1 512,944.29 sg13_lv_pmos
M$3111 \$2886 \$2887 \$2904 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $3112 r0 *1 516.84,944.265 sg13_lv_pmos
M$3112 VDD \$2896 \$2897 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3114 r0 *1 436.36,963.98 sg13_lv_pmos
M$3114 VDD \$2863 \$3053 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3115 r0 *1 437.44,963.825 sg13_lv_pmos
M$3115 \$3054 \$2897 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $3116 r0 *1 437.98,963.965 sg13_lv_pmos
M$3116 VDD \$2882 \$3055 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3117 r0 *1 438.49,963.965 sg13_lv_pmos
M$3117 \$3055 \$3054 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3118 r0 *1 439.93,964.105 sg13_lv_pmos
M$3118 VDD \$2882 \$3056 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $3119 r0 *1 440.44,964.105 sg13_lv_pmos
M$3119 VDD \$2897 \$3056 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $3120 r0 *1 440.95,963.965 sg13_lv_pmos
M$3120 VDD \$3056 \$3057 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3121 r0 *1 446.165,968.92 sg13_lv_pmos
M$3121 \$3093 \$3053 CORE$12 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $3124 r0 *1 448.83,969.565 sg13_lv_pmos
M$3124 \$3093 \$3055 PAD|VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $3125 r0 *1 454.21,968.655 sg13_lv_pmos
M$3125 \$3099 \$3099 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $3129 r0 *1 458.58,968.64 sg13_lv_pmos
M$3129 \$3048 \$3047 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $3133 r0 *1 465.44,963.98 sg13_lv_pmos
M$3133 VDD \$2882 \$3059 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3134 r0 *1 466.52,963.825 sg13_lv_pmos
M$3134 \$3060 \$2934 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $3135 r0 *1 467.06,963.965 sg13_lv_pmos
M$3135 VDD \$2863 \$3061 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3136 r0 *1 467.57,963.965 sg13_lv_pmos
M$3136 \$3061 \$3060 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3137 r0 *1 469.01,964.105 sg13_lv_pmos
M$3137 VDD \$2863 \$3062 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $3138 r0 *1 469.52,964.105 sg13_lv_pmos
M$3138 VDD \$2934 \$3062 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $3139 r0 *1 470.03,963.965 sg13_lv_pmos
M$3139 VDD \$3062 \$3063 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3140 r0 *1 475.245,968.92 sg13_lv_pmos
M$3140 \$3094 \$3059 \$3048 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $3143 r0 *1 477.91,969.565 sg13_lv_pmos
M$3143 \$3094 \$3061 PAD|VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $3144 r0 *1 483.29,968.655 sg13_lv_pmos
M$3144 \$3100 \$3100 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $3148 r0 *1 487.66,968.64 sg13_lv_pmos
M$3148 \$3050 \$3049 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $3152 r0 *1 515.9,949.25 sg13_lv_pmos
M$3152 VDD \$2897 \$3150 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3154 r0 *1 1056.005,997.48 sg13_lv_pmos
M$3154 \$3148 \$3150 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $3155 r0 *1 1056.005,1000.99 sg13_lv_pmos
M$3155 \$3176 \$3150 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $3156 r0 *1 700.255,1056.005 sg13_lv_pmos
M$3156 \$1474 \$3240 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $3157 r0 *1 800.255,1056.005 sg13_lv_pmos
M$3157 \$2651 \$3241 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $3158 r0 *1 900.255,1056.005 sg13_lv_pmos
M$3158 \$3013 \$3242 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $3159 r0 *1 501.765,243.945 sg13_hv_pmos
M$3159 VDD CORE \$178 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $3160 r0 *1 701.765,243.945 sg13_hv_pmos
M$3160 VDD CORE$1 \$179 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $3161 r0 *1 801.765,243.945 sg13_hv_pmos
M$3161 VDD CORE$2 \$180 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $3162 r0 *1 901.765,243.945 sg13_hv_pmos
M$3162 VDD CORE$3 \$181 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $3163 r0 *1 151.08,285.52 sg13_hv_pmos
M$3163 AVDD \$220 IN6|PAD AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3203 r0 *1 1141.82,294.58 sg13_hv_pmos
M$3203 IOVDD \$209 OUT6 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $3219 r0 *1 1068.82,297.64 sg13_hv_pmos
M$3219 \$231 \$241 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3220 r0 *1 1068.82,298.47 sg13_hv_pmos
M$3220 IOVDD \$231 \$241 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3221 r0 *1 1068.82,299.81 sg13_hv_pmos
M$3221 IOVDD \$241 \$249 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3222 r0 *1 1068.82,301.15 sg13_hv_pmos
M$3222 \$269 \$287 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3223 r0 *1 1068.82,301.98 sg13_hv_pmos
M$3223 IOVDD \$269 \$287 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3224 r0 *1 1068.82,303.32 sg13_hv_pmos
M$3224 IOVDD \$287 \$209 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3225 r0 *1 151.08,385.52 sg13_hv_pmos
M$3225 AVDD \$610 IN5|PAD AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3265 r0 *1 1141.82,394.58 sg13_hv_pmos
M$3265 IOVDD \$599 OUT5 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $3281 r0 *1 1068.82,397.64 sg13_hv_pmos
M$3281 \$644 \$665 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3282 r0 *1 1068.82,398.47 sg13_hv_pmos
M$3282 IOVDD \$644 \$665 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3283 r0 *1 1068.82,399.81 sg13_hv_pmos
M$3283 IOVDD \$665 \$672 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3284 r0 *1 1068.82,401.15 sg13_hv_pmos
M$3284 \$688 \$698 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3285 r0 *1 1068.82,401.98 sg13_hv_pmos
M$3285 IOVDD \$688 \$698 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3286 r0 *1 1068.82,403.32 sg13_hv_pmos
M$3286 IOVDD \$698 \$599 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3287 r0 *1 151.08,485.52 sg13_hv_pmos
M$3287 AVDD \$1074 IN4|PAD AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3327 r0 *1 1141.82,494.58 sg13_hv_pmos
M$3327 IOVDD \$1063 OUT4 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $3343 r0 *1 1068.82,497.64 sg13_hv_pmos
M$3343 \$1084 \$1097 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3344 r0 *1 1068.82,498.47 sg13_hv_pmos
M$3344 IOVDD \$1084 \$1097 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3345 r0 *1 1068.82,499.81 sg13_hv_pmos
M$3345 IOVDD \$1097 \$1100 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3346 r0 *1 1068.82,501.15 sg13_hv_pmos
M$3346 \$1112 \$1119 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3347 r0 *1 1068.82,501.98 sg13_hv_pmos
M$3347 IOVDD \$1112 \$1119 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3348 r0 *1 1068.82,503.32 sg13_hv_pmos
M$3348 IOVDD \$1119 \$1063 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3349 r0 *1 151.08,585.52 sg13_hv_pmos
M$3349 AVDD \$1467 PAD|VLO AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3389 r0 *1 151.08,685.52 sg13_hv_pmos
M$3389 AVDD \$1810 PAD|VHI AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3429 r0 *1 1125.09,678.44 sg13_hv_pmos
M$3429 IOVDD \$1802 \$1803 IOVDD sg13_hv_pmos W=350.0 L=0.5
* device instance $3479 r0 *1 151.08,785.52 sg13_hv_pmos
M$3479 AVDD \$1900 IN3|PAD AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3519 r0 *1 1141.82,794.58 sg13_hv_pmos
M$3519 IOVDD \$1889 OUT3 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $3535 r0 *1 1068.82,797.64 sg13_hv_pmos
M$3535 \$1910 \$1923 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3536 r0 *1 1068.82,798.47 sg13_hv_pmos
M$3536 IOVDD \$1910 \$1923 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3537 r0 *1 1068.82,799.81 sg13_hv_pmos
M$3537 IOVDD \$1923 \$1926 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3538 r0 *1 1068.82,801.15 sg13_hv_pmos
M$3538 \$1938 \$1945 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3539 r0 *1 1068.82,801.98 sg13_hv_pmos
M$3539 IOVDD \$1938 \$1945 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3540 r0 *1 1068.82,803.32 sg13_hv_pmos
M$3540 IOVDD \$1945 \$1889 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3541 r0 *1 531.375,828.1 sg13_hv_pmos
M$3541 IOVDD \$2126 PAD|VLDO IOVDD sg13_hv_pmos W=1414.0 L=0.44999999999999996
* device instance $3569 r0 *1 507.535,883.64 sg13_hv_pmos
M$3569 \$2545 \$2545 IOVDD IOVDD sg13_hv_pmos W=1.0 L=5.0
* device instance $3570 r0 *1 510.135,880.705 sg13_hv_pmos
M$3570 IOVDD \$2619 \$2619 IOVDD sg13_hv_pmos W=54.0 L=0.8999999999999999
* device instance $3588 r0 *1 539.845,885.93 sg13_hv_pmos
M$3588 IOVDD \$2560 \$2560 IOVDD sg13_hv_pmos W=36.0 L=0.8999999999999999
* device instance $3594 r0 *1 547.525,885.93 sg13_hv_pmos
M$3594 IOVDD \$2560 \$2126 IOVDD sg13_hv_pmos W=36.0 L=0.8999999999999999
* device instance $3600 r0 *1 158.18,885.52 sg13_hv_pmos
M$3600 AVDD \$2707 IN2|PAD AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3620 r0 *1 510.135,886.92 sg13_hv_pmos
M$3620 IOVDD \$2619 \$2544 IOVDD sg13_hv_pmos W=54.0 L=0.8999999999999999
* device instance $3658 r0 *1 1068.82,899.81 sg13_hv_pmos
M$3658 IOVDD \$2783 \$2789 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3659 r0 *1 1068.82,897.64 sg13_hv_pmos
M$3659 \$2774 \$2783 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3660 r0 *1 1068.82,898.47 sg13_hv_pmos
M$3660 IOVDD \$2774 \$2783 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3661 r0 *1 1141.82,894.58 sg13_hv_pmos
M$3661 IOVDD \$2683 OUT2 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $3677 r0 *1 1068.82,901.15 sg13_hv_pmos
M$3677 \$2801 \$2808 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3678 r0 *1 1068.82,901.98 sg13_hv_pmos
M$3678 IOVDD \$2801 \$2808 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3679 r0 *1 1068.82,903.32 sg13_hv_pmos
M$3679 IOVDD \$2808 \$2683 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3680 r0 *1 151.08,985.52 sg13_hv_pmos
M$3680 AVDD \$3139 IN1|PAD AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3720 r0 *1 1141.82,994.58 sg13_hv_pmos
M$3720 IOVDD \$3129 OUT1 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $3736 r0 *1 1068.82,997.64 sg13_hv_pmos
M$3736 \$3149 \$3159 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3737 r0 *1 1068.82,998.47 sg13_hv_pmos
M$3737 IOVDD \$3149 \$3159 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3738 r0 *1 1068.82,999.81 sg13_hv_pmos
M$3738 IOVDD \$3159 \$3165 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3739 r0 *1 1068.82,1001.15 sg13_hv_pmos
M$3739 \$3177 \$3184 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3740 r0 *1 1068.82,1001.98 sg13_hv_pmos
M$3740 IOVDD \$3177 \$3184 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3741 r0 *1 1068.82,1003.32 sg13_hv_pmos
M$3741 IOVDD \$3184 \$3129 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3742 r0 *1 701.765,1056.055 sg13_hv_pmos
M$3742 VDD CORE$13 \$3240 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $3743 r0 *1 801.765,1056.055 sg13_hv_pmos
M$3743 VDD CORE$14 \$3241 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $3744 r0 *1 901.765,1056.055 sg13_hv_pmos
M$3744 VDD CORE$15 \$3242 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $3745 r0 *1 278.44,1125.09 sg13_hv_pmos
M$3745 AVDD \$3368 \$3309 AVDD sg13_hv_pmos W=350.0 L=0.5
* device instance $3795 r0 *1 578.44,1125.09 sg13_hv_pmos
M$3795 IOVDD \$3369 \$3310 IOVDD sg13_hv_pmos W=350.0 L=0.5
* device instance $3845 r0 *1 978.44,1125.09 sg13_hv_pmos
M$3845 VDD \$3370 \$3311 VDD sg13_hv_pmos W=350.0 L=0.5
* device instance $3895 r0 *1 385.52,1148.92 sg13_hv_pmos
M$3895 AVDD \$3326 PAD|VREF AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3935 r0 *1 485.52,1148.92 sg13_hv_pmos
M$3935 AVDD \$3327 PAD|VLDO AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3975 r0 *1 264.54,104.19 dantenna
D$3975 VSS VSS dantenna A=35.0028 P=58.08 m=10
* device instance $3979 r0 *1 464.54,104.19 dantenna
D$3979 VSS PAD|RES dantenna A=35.0028 P=58.08 m=2
* device instance $3983 r0 *1 664.54,104.19 dantenna
D$3983 VSS CK4|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $3985 r0 *1 764.54,104.19 dantenna
D$3985 VSS CK5|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $3987 r0 *1 864.54,104.19 dantenna
D$3987 VSS CK6|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $3991 r0 *1 100.44,400 dantenna
D$3991 VSS IN5|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $3992 r0 *1 100.44,300 dantenna
D$3992 VSS IN6|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $3995 r0 *1 222.54,417.63 dantenna
D$3995 VSS CORE$5 dantenna A=1.984 P=7.48 m=1
* device instance $3996 r0 *1 222.54,317.63 dantenna
D$3996 VSS CORE$4 dantenna A=1.984 P=7.48 m=1
* device instance $3997 r0 *1 505.225,222.54 dantenna
D$3997 VSS CORE dantenna A=1.984 P=7.48 m=1
* device instance $3998 r0 *1 705.225,222.54 dantenna
D$3998 VSS CORE$1 dantenna A=1.984 P=7.48 m=1
* device instance $3999 r0 *1 805.225,222.54 dantenna
D$3999 VSS CORE$2 dantenna A=1.984 P=7.48 m=1
* device instance $4000 r0 *1 905.225,222.54 dantenna
D$4000 VSS CORE$3 dantenna A=1.984 P=7.48 m=1
* device instance $4001 r0 *1 1195.06,300 dantenna
D$4001 VSS OUT6 dantenna A=35.0028 P=58.08 m=2
* device instance $4002 r0 *1 1195.06,400 dantenna
D$4002 VSS OUT5 dantenna A=35.0028 P=58.08 m=2
* device instance $4005 r0 *1 1207.17,377.975 dantenna
D$4005 VSS \$672 dantenna A=0.192 P=1.88 m=1
* device instance $4006 r0 *1 1207.17,277.975 dantenna
D$4006 VSS \$249 dantenna A=0.192 P=1.88 m=1
* device instance $4007 r0 *1 1207.17,477.975 dantenna
D$4007 VSS \$1100 dantenna A=0.192 P=1.88 m=1
* device instance $4008 r0 *1 100.44,500 dantenna
D$4008 VSS IN4|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $4010 r0 *1 1195.06,500 dantenna
D$4010 VSS OUT4 dantenna A=35.0028 P=58.08 m=2
* device instance $4012 r0 *1 222.54,517.63 dantenna
D$4012 VSS CORE$6 dantenna A=1.984 P=7.48 m=1
* device instance $4015 r0 *1 100.44,600 dantenna
D$4015 VSS PAD|VLO dantenna A=35.0028 P=58.08 m=2
* device instance $4017 r0 *1 222.54,617.63 dantenna
D$4017 VSS CORE$7 dantenna A=1.984 P=7.48 m=1
* device instance $4018 r0 *1 1192.65,664.765 dantenna
D$4018 VSS \$1803 dantenna A=0.192 P=1.88 m=1
* device instance $4019 r0 *1 100.44,700 dantenna
D$4019 VSS PAD|VHI dantenna A=35.0028 P=58.08 m=2
* device instance $4021 r0 *1 222.54,717.63 dantenna
D$4021 VSS CORE$8 dantenna A=1.984 P=7.48 m=1
* device instance $4022 r0 *1 1207.17,777.975 dantenna
D$4022 VSS \$1926 dantenna A=0.192 P=1.88 m=1
* device instance $4023 r0 *1 100.44,800 dantenna
D$4023 VSS IN3|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $4025 r0 *1 1195.06,800 dantenna
D$4025 VSS OUT3 dantenna A=35.0028 P=58.08 m=2
* device instance $4027 r0 *1 222.54,817.63 dantenna
D$4027 VSS CORE$9 dantenna A=1.984 P=7.48 m=1
* device instance $4028 r0 *1 1207.17,877.975 dantenna
D$4028 VSS \$2789 dantenna A=0.192 P=1.88 m=1
* device instance $4029 r0 *1 100.44,900 dantenna
D$4029 VSS IN2|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $4031 r0 *1 1195.06,900 dantenna
D$4031 VSS OUT2 dantenna A=35.0028 P=58.08 m=2
* device instance $4033 r0 *1 222.54,917.63 dantenna
D$4033 VSS CORE$11 dantenna A=1.984 P=7.48 m=1
* device instance $4034 r0 *1 1207.17,977.975 dantenna
D$4034 VSS \$3165 dantenna A=0.192 P=1.88 m=1
* device instance $4035 r0 *1 100.44,1000 dantenna
D$4035 VSS IN1|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $4037 r0 *1 1195.06,1000 dantenna
D$4037 VSS OUT1 dantenna A=35.0028 P=58.08 m=2
* device instance $4039 r0 *1 222.54,1017.63 dantenna
D$4039 VSS CORE$12 dantenna A=1.984 P=7.48 m=1
* device instance $4040 r0 *1 417.63,1077.46 dantenna
D$4040 VSS CORE$10 dantenna A=1.984 P=7.48 m=1
* device instance $4041 r0 *1 517.63,1077.46 dantenna
D$4041 VSS CORE$16 dantenna A=1.984 P=7.48 m=1
* device instance $4042 r0 *1 705.225,1077.46 dantenna
D$4042 VSS CORE$13 dantenna A=1.984 P=7.48 m=1
* device instance $4043 r0 *1 805.225,1077.46 dantenna
D$4043 VSS CORE$14 dantenna A=1.984 P=7.48 m=1
* device instance $4044 r0 *1 905.225,1077.46 dantenna
D$4044 VSS CORE$15 dantenna A=1.984 P=7.48 m=1
* device instance $4045 r0 *1 664.54,1195.81 dantenna
D$4045 VSS CK3|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $4047 r0 *1 764.54,1195.81 dantenna
D$4047 VSS CK2|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $4049 r0 *1 864.54,1195.81 dantenna
D$4049 VSS CK1|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $4051 r0 *1 264.765,1192.65 dantenna
D$4051 VSS \$3309 dantenna A=0.192 P=1.88 m=1
* device instance $4052 r0 *1 400,1195.06 dantenna
D$4052 VSS PAD|VREF dantenna A=35.0028 P=58.08 m=2
* device instance $4053 r0 *1 500,1195.06 dantenna
D$4053 VSS PAD|VLDO dantenna A=35.0028 P=58.08 m=2
* device instance $4054 r0 *1 564.765,1192.65 dantenna
D$4054 VSS \$3310 dantenna A=0.192 P=1.88 m=1
* device instance $4055 r0 *1 964.765,1192.65 dantenna
D$4055 VSS \$3311 dantenna A=0.192 P=1.88 m=1
* device instance $4058 r0 *1 264.54,163.19 dpantenna
D$4058 VSS AVDD dpantenna A=35.0028 P=58.08 m=4
* device instance $4062 r0 *1 464.54,163.19 dpantenna
D$4062 PAD|RES IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4064 r0 *1 564.54,163.19 dpantenna
D$4064 VSS IOVDD dpantenna A=35.0028 P=58.08 m=6
* device instance $4066 r0 *1 664.54,163.19 dpantenna
D$4066 CK4|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4068 r0 *1 764.54,163.19 dpantenna
D$4068 CK5|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4070 r0 *1 864.54,163.19 dpantenna
D$4070 CK6|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4074 r0 *1 227.51,315.46 dpantenna
D$4074 CORE$4 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4075 r0 *1 227.51,415.46 dpantenna
D$4075 CORE$5 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4076 r0 *1 227.51,515.46 dpantenna
D$4076 CORE$6 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4077 r0 *1 227.51,615.46 dpantenna
D$4077 CORE$7 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4078 r0 *1 227.51,715.46 dpantenna
D$4078 CORE$8 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4079 r0 *1 227.51,815.46 dpantenna
D$4079 CORE$9 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4080 r0 *1 227.51,915.46 dpantenna
D$4080 CORE$11 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4081 r0 *1 227.51,1015.46 dpantenna
D$4081 CORE$12 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4082 r0 *1 415.46,1072.49 dpantenna
D$4082 CORE$10 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4083 r0 *1 515.46,1072.49 dpantenna
D$4083 CORE$16 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4084 r0 *1 503.055,227.51 dpantenna
D$4084 CORE IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4085 r0 *1 703.055,227.51 dpantenna
D$4085 CORE$1 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4086 r0 *1 803.055,227.51 dpantenna
D$4086 CORE$2 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4087 r0 *1 903.055,227.51 dpantenna
D$4087 CORE$3 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4088 r0 *1 703.055,1072.49 dpantenna
D$4088 CORE$13 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4089 r0 *1 803.055,1072.49 dpantenna
D$4089 CORE$14 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4090 r0 *1 903.055,1072.49 dpantenna
D$4090 CORE$15 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4091 r0 *1 1138.81,277.975 dpantenna
D$4091 \$209 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $4092 r0 *1 135.96,300 dpantenna
D$4092 IN6|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4094 r0 *1 1159.54,300 dpantenna
D$4094 OUT6 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4096 r0 *1 135.96,400 dpantenna
D$4096 IN5|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4098 r0 *1 1138.81,377.975 dpantenna
D$4098 \$599 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $4099 r0 *1 1159.54,400 dpantenna
D$4099 OUT5 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4101 r0 *1 135.96,500 dpantenna
D$4101 IN4|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4103 r0 *1 1138.81,477.975 dpantenna
D$4103 \$1063 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $4104 r0 *1 1159.54,500 dpantenna
D$4104 OUT4 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4106 r0 *1 135.96,600 dpantenna
D$4106 PAD|VLO AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4110 r0 *1 135.96,700 dpantenna
D$4110 PAD|VHI AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4112 r0 *1 1138.81,777.975 dpantenna
D$4112 \$1889 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $4113 r0 *1 135.96,800 dpantenna
D$4113 IN3|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4115 r0 *1 1159.54,800 dpantenna
D$4115 OUT3 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4117 r0 *1 135.96,900 dpantenna
D$4117 IN2|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4119 r0 *1 1138.81,877.975 dpantenna
D$4119 \$2683 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $4120 r0 *1 1159.54,900 dpantenna
D$4120 OUT2 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4122 r0 *1 135.96,1000 dpantenna
D$4122 IN1|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4124 r0 *1 1138.81,977.975 dpantenna
D$4124 \$3129 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $4125 r0 *1 1159.54,1000 dpantenna
D$4125 OUT1 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4127 r0 *1 664.54,1136.81 dpantenna
D$4127 CK3|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4129 r0 *1 764.54,1136.81 dpantenna
D$4129 CK2|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4131 r0 *1 864.54,1136.81 dpantenna
D$4131 CK1|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4133 r0 *1 400,1159.54 dpantenna
D$4133 PAD|VREF AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4135 r0 *1 500,1159.54 dpantenna
D$4135 PAD|VLDO AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4137 r0 *1 500.685,221.11 rppd
R$4137 PAD|RES CORE rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4138 r0 *1 700.685,221.11 rppd
R$4138 CK4|PAD CORE$1 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4139 r0 *1 800.685,221.11 rppd
R$4139 CK5|PAD CORE$2 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4140 r0 *1 900.685,221.11 rppd
R$4140 CK6|PAD CORE$3 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4141 r0 *1 88.75,326.305 rppd
R$4141 VSS \$219 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4142 r0 *1 147.75,326.305 rppd
R$4142 AVDD \$220 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4143 r0 *1 221.11,313.09 rppd
R$4143 IN6|PAD CORE$4 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4144 r0 *1 88.75,426.305 rppd
R$4144 VSS \$609 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4145 r0 *1 147.75,426.305 rppd
R$4145 AVDD \$610 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4146 r0 *1 221.11,413.09 rppd
R$4146 IN5|PAD CORE$5 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4147 r0 *1 88.75,526.305 rppd
R$4147 VSS \$1073 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4148 r0 *1 147.75,526.305 rppd
R$4148 AVDD \$1074 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4149 r0 *1 221.11,513.09 rppd
R$4149 IN4|PAD CORE$6 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4150 r0 *1 88.75,626.305 rppd
R$4150 VSS \$1466 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4151 r0 *1 147.75,626.305 rppd
R$4151 AVDD \$1467 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4152 r0 *1 221.11,613.09 rppd
R$4152 PAD|VLO CORE$7 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4153 r0 *1 1161.29,678.875 rppd
R$4153 IOVDD \$1802 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $4154 r0 *1 221.11,713.09 rppd
R$4154 PAD|VHI CORE$8 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4155 r0 *1 88.75,726.305 rppd
R$4155 VSS \$1809 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4156 r0 *1 147.75,726.305 rppd
R$4156 AVDD \$1810 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4157 r0 *1 88.75,826.305 rppd
R$4157 VSS \$1899 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4158 r0 *1 147.75,826.305 rppd
R$4158 AVDD \$1900 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4159 r0 *1 221.11,813.09 rppd
R$4159 IN3|PAD CORE$9 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4160 r0 *1 221.11,913.09 rppd
R$4160 IN2|PAD CORE$11 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4161 r0 *1 88.75,926.305 rppd
R$4161 VSS \$2706 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4162 r0 *1 147.75,926.305 rppd
R$4162 AVDD \$2707 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4163 r0 *1 88.75,1026.305 rppd
R$4163 VSS \$3138 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4164 r0 *1 147.75,1026.305 rppd
R$4164 AVDD \$3139 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4165 r0 *1 221.11,1013.09 rppd
R$4165 IN1|PAD CORE$12 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4166 r0 *1 413.09,1076.03 rppd
R$4166 CORE$10 PAD|VREF rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4167 r0 *1 513.09,1076.03 rppd
R$4167 CORE$16 PAD|VLDO rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4168 r0 *1 700.685,1076.03 rppd
R$4168 CORE$13 CK3|PAD rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4169 r0 *1 800.685,1076.03 rppd
R$4169 CORE$14 CK2|PAD rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4170 r0 *1 900.685,1076.03 rppd
R$4170 CORE$15 CK1|PAD rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4171 r0 *1 278.875,1161.29 rppd
R$4171 AVDD \$3368 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $4172 r0 *1 426.305,1138.49 rppd
R$4172 \$3326 AVDD rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4173 r0 *1 526.305,1138.49 rppd
R$4173 \$3327 AVDD rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4174 r0 *1 578.875,1161.29 rppd
R$4174 IOVDD \$3369 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $4175 r0 *1 978.875,1161.29 rppd
R$4175 VDD \$3370 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $4176 r0 *1 426.305,1206.85 rppd
R$4176 \$3440 VSS rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4177 r0 *1 526.305,1206.85 rppd
R$4177 \$3441 VSS rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4178 r0 *1 518.845,859.565 rhigh
R$4178 VSS \$2592 rhigh w=0.5 l=0.96 ps=0 b=0 m=2
* device instance $4180 r0 *1 555.805,883.57 rhigh
R$4180 \$2126 \$2129 rhigh w=0.5 l=3.84 ps=0 b=0 m=1
* device instance $4184 r0 *1 463.265,300.165 cap_cmim
C$4184 \$272 \$248 cap_cmim w=8.16 l=8.16 m=1
* device instance $4185 r0 *1 463.27,309.855 cap_cmim
C$4185 \$298 \$271 cap_cmim w=8.16 l=8.16 m=1
* device instance $4186 r0 *1 455.04,311.655 cap_cmim
C$4186 \$248 \$347 cap_cmim w=5.77 l=5.77 m=1
* device instance $4187 r0 *1 438.16,318.59 cap_cmim
C$4187 \$440 \$437 cap_cmim w=8.16 l=8.16 m=1
* device instance $4188 r0 *1 438.165,328.28 cap_cmim
C$4188 \$449 \$346 cap_cmim w=8.16 l=8.16 m=1
* device instance $4189 r0 *1 429.935,330.08 cap_cmim
C$4189 \$437 \$480 cap_cmim w=5.77 l=5.77 m=1
* device instance $4190 r0 *1 439.895,391.265 cap_cmim
C$4190 \$615 \$616 cap_cmim w=8.16 l=8.16 m=1
* device instance $4191 r0 *1 449.03,330.495 cap_cmim
C$4191 \$526 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $4192 r0 *1 492.37,391.265 cap_cmim
C$4192 \$618 \$617 cap_cmim w=8.16 l=8.16 m=1
* device instance $4193 r0 *1 449.47,391.27 cap_cmim
C$4193 \$616 \$632 cap_cmim w=5.77 l=5.77 m=1
* device instance $4194 r0 *1 457.715,410.955 cap_cmim
C$4194 \$754 \$799 cap_cmim w=8.16 l=8.16 m=1
* device instance $4195 r0 *1 474.55,410.955 cap_cmim
C$4195 \$755 \$795 cap_cmim w=8.16 l=8.16 m=1
* device instance $4196 r0 *1 485.185,391.27 cap_cmim
C$4196 \$617 \$659 cap_cmim w=5.77 l=5.77 m=1
* device instance $4197 r0 *1 471.465,445.3 cap_cmim
C$4197 \$961 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $4198 r0 *1 473.165,512.175 cap_cmim
C$4198 \$1183 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $4199 r0 *1 430.955,540.41 cap_cmim
C$4199 \$1412 \$1401 cap_cmim w=5.77 l=5.77 m=1
* device instance $4200 r0 *1 465.955,540.41 cap_cmim
C$4200 \$1413 \$1402 cap_cmim w=5.77 l=5.77 m=1
* device instance $4201 r0 *1 439.56,542.23 cap_cmim
C$4201 \$1377 \$1412 cap_cmim w=8.16 l=8.16 m=1
* device instance $4202 r0 *1 474.56,542.23 cap_cmim
C$4202 \$1378 \$1413 cap_cmim w=8.16 l=8.16 m=1
* device instance $4203 r0 *1 443.88,615.55 cap_cmim
C$4203 \$1612 \$1653 cap_cmim w=5.77 l=5.77 m=1
* device instance $4204 r0 *1 450.88,542.235 cap_cmim
C$4204 \$1372 \$1414 cap_cmim w=8.16 l=8.16 m=1
* device instance $4205 r0 *1 479.935,615.55 cap_cmim
C$4205 \$1613 \$1654 cap_cmim w=5.77 l=5.77 m=1
* device instance $4206 r0 *1 485.88,542.235 cap_cmim
C$4206 \$1182 \$1411 cap_cmim w=8.16 l=8.16 m=1
* device instance $4207 r0 *1 509.38,615.465 cap_cmim
C$4207 \$1679 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $4208 r0 *1 430.19,624.19 cap_cmim
C$4208 \$1689 \$1633 cap_cmim w=8.16 l=8.16 m=1
* device instance $4209 r0 *1 466.245,624.19 cap_cmim
C$4209 \$1690 \$1634 cap_cmim w=8.16 l=8.16 m=1
* device instance $4210 r0 *1 441.11,625.165 cap_cmim
C$4210 \$1723 \$1612 cap_cmim w=8.16 l=8.16 m=1
* device instance $4211 r0 *1 477.165,625.165 cap_cmim
C$4211 \$1724 \$1613 cap_cmim w=8.16 l=8.16 m=1
* device instance $4212 r0 *1 429.41,680.555 cap_cmim
C$4212 VSS PAD|VLDO cap_cmim w=70 l=75 m=6
* device instance $4218 r0 *1 429.41,826.865 cap_cmim
C$4218 \$2129 PAD|VLDO cap_cmim w=60 l=60 m=1
* device instance $4219 r0 *1 623.755,834.77 cap_cmim
C$4219 \$2174 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $4220 r0 *1 576.305,835.415 cap_cmim
C$4220 \$2180 \$2261 cap_cmim w=8.16 l=8.16 m=1
* device instance $4221 r0 *1 587.54,835.275 cap_cmim
C$4221 \$2172 \$2164 cap_cmim w=8.16 l=8.16 m=1
* device instance $4222 r0 *1 597.895,835.415 cap_cmim
C$4222 \$2181 \$2262 cap_cmim w=8.16 l=8.16 m=1
* device instance $4223 r0 *1 609.13,835.275 cap_cmim
C$4223 \$2173 \$2209 cap_cmim w=8.16 l=8.16 m=1
* device instance $4224 r0 *1 576.185,848.635 cap_cmim
C$4224 \$2261 \$2256 cap_cmim w=5.77 l=5.77 m=1
* device instance $4225 r0 *1 597.775,848.635 cap_cmim
C$4225 \$2262 \$2257 cap_cmim w=5.77 l=5.77 m=1
* device instance $4226 r0 *1 484.5,930.31 cap_cmim
C$4226 \$2861 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $4227 r0 *1 435.61,966.96 cap_cmim
C$4227 \$3058 \$3093 cap_cmim w=5.77 l=5.77 m=1
* device instance $4228 r0 *1 464.69,966.96 cap_cmim
C$4228 \$3064 \$3094 cap_cmim w=5.77 l=5.77 m=1
* device instance $4229 r0 *1 434.36,974.655 cap_cmim
C$4229 \$3047 \$3058 cap_cmim w=8.16 l=8.16 m=1
* device instance $4230 r0 *1 463.44,974.655 cap_cmim
C$4230 \$3049 \$3064 cap_cmim w=8.16 l=8.16 m=1
* device instance $4231 r0 *1 450.71,975.895 cap_cmim
C$4231 \$3046 \$3048 cap_cmim w=8.16 l=8.16 m=1
* device instance $4232 r0 *1 479.79,975.895 cap_cmim
C$4232 \$3065 \$3050 cap_cmim w=8.16 l=8.16 m=1
.ENDS UHEE628_S2024

* Extracted by KLayout with SG13G2 LVS runset on : 02/05/2024 06:12

* cell sg13g2_RCClampInverter
.SUBCKT sg13g2_RCClampInverter
* device instance $1 r0 *1 7.72,6.54 sg13_hv_nmos
M$1 sub!$1 \$3 sub!$1 sub!$1 sg13_hv_nmos W=125.99999999999999
+ L=9.499999999999996
* device instance $8 r0 *1 72.38,6.54 sg13_hv_nmos
M$8 sub!$1 \$3 \$5 sub!$1 sg13_hv_nmos W=107.99999999999999 L=0.4999999999999999
* device instance $27 r0 *1 18.44,29.91 sg13_hv_pmos
M$27 \$8 \$3 \$5 \$8 sg13_hv_pmos W=349.99999999999994 L=0.4999999999999999
.ENDS sg13g2_RCClampInverter

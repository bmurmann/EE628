* Extracted by KLayout with SG13G2 LVS runset on : 04/05/2024 04:48

* cell IDSM2_T4
* pin sub!
.SUBCKT IDSM2_T4 sub!
* device instance $1 r0 *1 55.618,1.632 sg13_lv_nmos
M$1 \$14 \$11 \$24 sub! sg13_lv_nmos W=0.41999999999999993 L=0.12999999999999995
* device instance $2 r0 *1 56.008,1.632 sg13_lv_nmos
M$2 \$24 \$15 sub! sub! sg13_lv_nmos W=0.41999999999999993 L=0.12999999999999995
* device instance $3 r0 *1 56.568,1.632 sg13_lv_nmos
M$3 sub! \$2 \$25 sub! sg13_lv_nmos W=0.41999999999999993 L=0.12999999999999995
* device instance $4 r0 *1 56.923,1.632 sg13_lv_nmos
M$4 \$25 \$14 \$15 sub! sg13_lv_nmos W=0.41999999999999993 L=0.12999999999999995
* device instance $5 r0 *1 53.978,1.742 sg13_lv_nmos
M$5 sub! \$12 \$13 sub! sg13_lv_nmos W=0.6399999999999999 L=0.12999999999999995
* device instance $6 r0 *1 54.648,1.742 sg13_lv_nmos
M$6 \$13 \$3 \$14 sub! sg13_lv_nmos W=0.6399999999999999 L=0.12999999999999995
* device instance $7 r0 *1 52.098,1.857 sg13_lv_nmos
M$7 \$10 \$11 \$12 sub! sg13_lv_nmos W=0.41999999999999993 L=0.12999999999999995
* device instance $8 r0 *1 52.608,1.857 sg13_lv_nmos
M$8 \$12 \$3 \$23 sub! sg13_lv_nmos W=0.41999999999999993 L=0.12999999999999995
* device instance $9 r0 *1 52.998,1.857 sg13_lv_nmos
M$9 \$23 \$13 \$22 sub! sg13_lv_nmos W=0.41999999999999993 L=0.12999999999999995
* device instance $10 r0 *1 53.358,1.857 sg13_lv_nmos
M$10 sub! \$2 \$22 sub! sg13_lv_nmos W=0.41999999999999993 L=0.12999999999999995
* device instance $11 r0 *1 46.768,1.797 sg13_lv_nmos
M$11 sub! \$150 \$9 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $12 r0 *1 57.963,1.797 sg13_lv_nmos
M$12 sub! \$14 \$16 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $13 r0 *1 59.163,1.702 sg13_lv_nmos
M$13 \$17 \$14 sub! sub! sg13_lv_nmos W=0.5499999999999999 L=0.12999999999999995
* device instance $14 r0 *1 59.703,1.797 sg13_lv_nmos
M$14 sub! \$17 \$36 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $15 r0 *1 61.898,1.797 sg13_lv_nmos
M$15 sub! \$36 \$18 sub! sg13_lv_nmos W=1.4799999999999998 L=0.12999999999999995
* device instance $17 r0 *1 64.693,1.796 sg13_lv_nmos
M$17 sub! \$26 \$2 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $18 r0 *1 66.608,1.796 sg13_lv_nmos
M$18 sub! \$27 \$19 sub! sg13_lv_nmos W=1.4799999999999998 L=0.12999999999999995
* device instance $20 r0 *1 67.628,1.846 sg13_lv_nmos
M$20 sub! \$68 \$27 sub! sg13_lv_nmos W=0.6399999999999999 L=0.12999999999999995
* device instance $21 r0 *1 48.818,1.657 sg13_lv_nmos
M$21 \$10 \$68 \$21 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $22 r0 *1 49.188,1.657 sg13_lv_nmos
M$22 \$21 \$2 sub! sub! sg13_lv_nmos W=0.41999999999999993 L=0.12999999999999995
* device instance $23 r0 *1 50.333,1.972 sg13_lv_nmos
M$23 sub! \$150 \$11 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $24 r0 *1 50.843,1.972 sg13_lv_nmos
M$24 sub! \$11 \$3 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $25 r0 *1 51.503,8.202 sg13_lv_nmos
M$25 sub! \$58 \$59 sub! sg13_lv_nmos W=1.9999999999999996 L=0.9999999999999998
* device instance $26 r0 *1 51.703,10.304 sg13_lv_nmos
M$26 \$59 \$95 \$63 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $27 r0 *1 53.503,6.672 sg13_lv_nmos
M$27 \$48 \$150 \$49 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $28 r0 *1 52.903,10.304 sg13_lv_nmos
M$28 \$63 \$74 \$64 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $29 r0 *1 54.103,10.304 sg13_lv_nmos
M$29 \$74 \$64 \$65 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $30 r0 *1 55.503,8.202 sg13_lv_nmos
M$30 sub! \$49 \$60 sub! sg13_lv_nmos W=1.9999999999999996 L=0.9999999999999998
* device instance $31 r0 *1 55.303,10.304 sg13_lv_nmos
M$31 \$65 \$95 \$60 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $32 r0 *1 58.561,10.304 sg13_lv_nmos
M$32 sub! \$74 \$66 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $33 r0 *1 59.761,10.304 sg13_lv_nmos
M$33 \$66 \$68 \$67 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $34 r0 *1 60.961,10.304 sg13_lv_nmos
M$34 \$68 \$67 \$69 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $35 r0 *1 62.161,10.304 sg13_lv_nmos
M$35 \$69 \$64 sub! sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $36 r0 *1 8.155,16.051 sg13_lv_nmos
M$36 sub! \$86 \$87 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $40 r0 *1 11.035,16.051 sg13_lv_nmos
M$40 sub! \$87 \$88 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $44 r0 *1 13.915,16.051 sg13_lv_nmos
M$44 sub! \$88 \$89 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $48 r0 *1 16.795,16.051 sg13_lv_nmos
M$48 sub! \$89 \$90 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $52 r0 *1 19.675,16.051 sg13_lv_nmos
M$52 sub! \$90 \$91 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $56 r0 *1 22.555,16.051 sg13_lv_nmos
M$56 sub! \$91 \$92 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $60 r0 *1 28.315,16.051 sg13_lv_nmos
M$60 sub! \$93 \$94 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $64 r0 *1 31.135,16.051 sg13_lv_nmos
M$64 sub! \$94 \$95 sub! sg13_lv_nmos W=5.92 L=0.12999999999999995
* device instance $72 r0 *1 1.455,18.486 sg13_lv_nmos
M$72 sub! \$137 \$96 sub! sg13_lv_nmos W=1.4799999999999998
+ L=0.12999999999999995
* device instance $74 r0 *1 3.375,18.486 sg13_lv_nmos
M$74 sub! \$96 \$138 sub! sg13_lv_nmos W=1.4799999999999998
+ L=0.12999999999999995
* device instance $76 r0 *1 5.35,18.461 sg13_lv_nmos
M$76 \$139 \$92 sub! sub! sg13_lv_nmos W=1.4399999999999997
+ L=0.12999999999999998
* device instance $78 r0 *1 6.38,18.461 sg13_lv_nmos
M$78 \$139 \$138 \$140 sub! sg13_lv_nmos W=1.4399999999999997
+ L=0.12999999999999998
* device instance $80 r0 *1 5.35,16.076 sg13_lv_nmos
M$80 \$107 \$146 sub! sub! sg13_lv_nmos W=1.4399999999999997
+ L=0.12999999999999998
* device instance $82 r0 *1 6.38,16.076 sg13_lv_nmos
M$82 \$107 \$96 \$86 sub! sg13_lv_nmos W=1.4399999999999997
+ L=0.12999999999999998
* device instance $84 r0 *1 8.155,18.486 sg13_lv_nmos
M$84 sub! \$140 \$141 sub! sg13_lv_nmos W=2.9599999999999995
+ L=0.12999999999999995
* device instance $88 r0 *1 11.035,18.486 sg13_lv_nmos
M$88 sub! \$141 \$142 sub! sg13_lv_nmos W=2.9599999999999995
+ L=0.12999999999999995
* device instance $92 r0 *1 13.915,18.486 sg13_lv_nmos
M$92 sub! \$142 \$143 sub! sg13_lv_nmos W=2.9599999999999995
+ L=0.12999999999999995
* device instance $96 r0 *1 16.795,18.486 sg13_lv_nmos
M$96 sub! \$143 \$144 sub! sg13_lv_nmos W=2.9599999999999995
+ L=0.12999999999999995
* device instance $100 r0 *1 19.675,18.486 sg13_lv_nmos
M$100 sub! \$144 \$145 sub! sg13_lv_nmos W=2.9599999999999995
+ L=0.12999999999999995
* device instance $104 r0 *1 22.555,18.486 sg13_lv_nmos
M$104 sub! \$145 \$146 sub! sg13_lv_nmos W=2.9599999999999995
+ L=0.12999999999999995
* device instance $108 r0 *1 25.51,16.076 sg13_lv_nmos
M$108 \$108 \$92 sub! sub! sg13_lv_nmos W=1.4399999999999997
+ L=0.12999999999999998
* device instance $110 r0 *1 26.54,16.076 sg13_lv_nmos
M$110 \$108 \$90 \$93 sub! sg13_lv_nmos W=1.4399999999999997
+ L=0.12999999999999998
* device instance $112 r0 *1 25.51,18.461 sg13_lv_nmos
M$112 \$147 \$146 sub! sub! sg13_lv_nmos W=1.4399999999999997
+ L=0.12999999999999998
* device instance $114 r0 *1 26.54,18.461 sg13_lv_nmos
M$114 \$147 \$144 \$148 sub! sg13_lv_nmos W=1.4399999999999997
+ L=0.12999999999999998
* device instance $116 r0 *1 28.315,18.486 sg13_lv_nmos
M$116 sub! \$148 \$149 sub! sg13_lv_nmos W=2.9599999999999995
+ L=0.12999999999999995
* device instance $120 r0 *1 31.135,18.486 sg13_lv_nmos
M$120 sub! \$149 \$150 sub! sg13_lv_nmos W=5.92 L=0.12999999999999995
* device instance $128 r0 *1 1.5,32.466 sg13_lv_nmos
M$128 sub! \$150 \$186 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $129 r0 *1 2.935,32.561 sg13_lv_nmos
M$129 sub! \$36 \$187 sub! sg13_lv_nmos W=0.5499999999999999
+ L=0.12999999999999995
* device instance $130 r0 *1 3.785,32.466 sg13_lv_nmos
M$130 sub! \$95 \$200 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $131 r0 *1 4.095,32.466 sg13_lv_nmos
M$131 \$200 \$187 \$188 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $132 r0 *1 4.07,50.411 sg13_lv_nmos
M$132 \$235 \$190 \$263 sub! sg13_lv_nmos W=0.4999999999999999
+ L=0.12999999999999998
* device instance $133 r0 *1 5.785,32.626 sg13_lv_nmos
M$133 \$189 \$95 \$202 sub! sg13_lv_nmos W=0.6399999999999999
+ L=0.12999999999999995
* device instance $134 r0 *1 6.295,32.626 sg13_lv_nmos
M$134 sub! \$36 \$202 sub! sg13_lv_nmos W=0.6399999999999999
+ L=0.12999999999999995
* device instance $135 r0 *1 6.805,32.576 sg13_lv_nmos
M$135 sub! \$189 \$190 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $136 r0 *1 6.815,50.421 sg13_lv_nmos
M$136 \$235 \$150 \$248 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $137 r0 *1 13.55,32.481 sg13_lv_nmos
M$137 sub! \$191 \$191 sub! sg13_lv_nmos W=2.4999999999999996
+ L=1.4999999999999996
* device instance $138 r0 *1 14.09,50.376 sg13_lv_nmos
M$138 \$191 \$145 \$236 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $139 r0 *1 25.2,32.466 sg13_lv_nmos
M$139 sub! \$212 \$197 sub! sg13_lv_nmos W=2.4999999999999996
+ L=1.4999999999999996
* device instance $140 r0 *1 24.14,50.371 sg13_lv_nmos
M$140 \$236 \$95 \$247 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $141 r0 *1 25.45,50.371 sg13_lv_nmos
M$141 \$247 \$150 \$212 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $142 r0 *1 26.763,50.371 sg13_lv_nmos
M$142 \$247 \$26 \$197 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $143 r0 *1 36.5,32.466 sg13_lv_nmos
M$143 sub! \$95 \$192 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $144 r0 *1 37.935,32.561 sg13_lv_nmos
M$144 sub! \$19 \$193 sub! sg13_lv_nmos W=0.5499999999999999
+ L=0.12999999999999995
* device instance $145 r0 *1 38.785,32.466 sg13_lv_nmos
M$145 sub! \$150 \$211 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $146 r0 *1 39.095,32.466 sg13_lv_nmos
M$146 \$211 \$193 \$194 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $147 r0 *1 39.07,50.411 sg13_lv_nmos
M$147 \$249 \$196 \$263 sub! sg13_lv_nmos W=0.4999999999999999
+ L=0.12999999999999998
* device instance $148 r0 *1 40.785,32.626 sg13_lv_nmos
M$148 \$195 \$150 \$209 sub! sg13_lv_nmos W=0.6399999999999999
+ L=0.12999999999999995
* device instance $149 r0 *1 41.295,32.626 sg13_lv_nmos
M$149 sub! \$19 \$209 sub! sg13_lv_nmos W=0.6399999999999999
+ L=0.12999999999999995
* device instance $150 r0 *1 41.805,32.576 sg13_lv_nmos
M$150 sub! \$195 \$196 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $151 r0 *1 41.815,50.421 sg13_lv_nmos
M$151 \$249 \$95 \$197 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $152 r0 *1 48.55,32.481 sg13_lv_nmos
M$152 sub! \$58 \$58 sub! sg13_lv_nmos W=2.4999999999999996 L=1.4999999999999996
* device instance $153 r0 *1 49.09,50.376 sg13_lv_nmos
M$153 \$58 \$91 \$246 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $154 r0 *1 60.2,32.466 sg13_lv_nmos
M$154 sub! \$213 \$48 sub! sg13_lv_nmos W=2.4999999999999996
+ L=1.4999999999999996
* device instance $155 r0 *1 59.14,50.371 sg13_lv_nmos
M$155 \$246 \$150 \$237 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $156 r0 *1 60.45,50.371 sg13_lv_nmos
M$156 \$237 \$95 \$213 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $157 r0 *1 61.763,50.371 sg13_lv_nmos
M$157 \$237 \$26 \$48 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $158 r0 *1 54.613,3.292 sg13_lv_pmos
M$158 \$83 \$12 \$13 \$83 sg13_lv_pmos W=0.9999999999999998
+ L=0.12999999999999998
* device instance $159 r0 *1 55.123,3.292 sg13_lv_pmos
M$159 \$13 \$11 \$14 \$83 sg13_lv_pmos W=0.9999999999999998
+ L=0.12999999999999998
* device instance $160 r0 *1 55.773,3.622 sg13_lv_pmos
M$160 \$14 \$3 \$45 \$83 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $161 r0 *1 56.108,3.622 sg13_lv_pmos
M$161 \$45 \$15 \$83 \$83 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $162 r0 *1 56.618,3.622 sg13_lv_pmos
M$162 \$83 \$2 \$15 \$83 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $163 r0 *1 57.128,3.622 sg13_lv_pmos
M$163 \$83 \$14 \$15 \$83 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $164 r0 *1 57.688,3.457 sg13_lv_pmos
M$164 \$83 \$14 \$16 \$83 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $165 r0 *1 67.628,3.471 sg13_lv_pmos
M$165 \$83 \$68 \$27 \$83 sg13_lv_pmos W=0.9999999999999998
+ L=0.12999999999999998
* device instance $166 r0 *1 66.608,3.456 sg13_lv_pmos
M$166 \$83 \$27 \$19 \$83 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $168 r0 *1 59.163,3.597 sg13_lv_pmos
M$168 \$83 \$14 \$17 \$83 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $169 r0 *1 59.673,3.457 sg13_lv_pmos
M$169 \$83 \$17 \$36 \$83 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $170 r0 *1 61.888,3.457 sg13_lv_pmos
M$170 \$83 \$36 \$18 \$83 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $172 r0 *1 46.778,3.472 sg13_lv_pmos
M$172 \$83 \$150 \$9 \$83 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $173 r0 *1 50.303,3.517 sg13_lv_pmos
M$173 \$11 \$150 \$83 \$83 sg13_lv_pmos W=0.9999999999999998
+ L=0.12999999999999998
* device instance $174 r0 *1 50.813,3.517 sg13_lv_pmos
M$174 \$83 \$11 \$3 \$83 sg13_lv_pmos W=0.9999999999999998 L=0.12999999999999998
* device instance $175 r0 *1 51.973,3.582 sg13_lv_pmos
M$175 \$10 \$3 \$12 \$83 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $176 r0 *1 52.483,3.582 sg13_lv_pmos
M$176 \$12 \$11 \$41 \$83 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $177 r0 *1 52.858,3.582 sg13_lv_pmos
M$177 \$41 \$13 \$83 \$83 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $178 r0 *1 53.433,3.582 sg13_lv_pmos
M$178 \$83 \$2 \$12 \$83 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $179 r0 *1 64.703,3.471 sg13_lv_pmos
M$179 \$83 \$26 \$2 \$83 sg13_lv_pmos W=1.1199999999999999 L=0.12999999999999995
* device instance $180 r0 *1 5.35,14.391 sg13_lv_pmos
M$180 \$83 \$146 \$86 \$83 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $182 r0 *1 6.38,14.391 sg13_lv_pmos
M$182 \$83 \$96 \$86 \$83 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $184 r0 *1 8.155,14.391 sg13_lv_pmos
M$184 \$83 \$86 \$87 \$83 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $188 r0 *1 11.035,14.391 sg13_lv_pmos
M$188 \$83 \$87 \$88 \$83 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $192 r0 *1 13.915,14.391 sg13_lv_pmos
M$192 \$83 \$88 \$89 \$83 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $196 r0 *1 16.795,14.391 sg13_lv_pmos
M$196 \$83 \$89 \$90 \$83 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $200 r0 *1 19.675,14.391 sg13_lv_pmos
M$200 \$83 \$90 \$91 \$83 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $204 r0 *1 22.555,14.391 sg13_lv_pmos
M$204 \$83 \$91 \$92 \$83 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $208 r0 *1 25.51,14.391 sg13_lv_pmos
M$208 \$83 \$92 \$93 \$83 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $210 r0 *1 26.54,14.391 sg13_lv_pmos
M$210 \$83 \$90 \$93 \$83 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $212 r0 *1 28.315,14.391 sg13_lv_pmos
M$212 \$83 \$93 \$94 \$83 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $216 r0 *1 31.135,14.391 sg13_lv_pmos
M$216 \$83 \$94 \$95 \$83 sg13_lv_pmos W=8.959999999999999 L=0.12999999999999995
* device instance $224 r0 *1 48.773,3.807 sg13_lv_pmos
M$224 \$83 \$68 \$10 \$83 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $225 r0 *1 49.283,3.807 sg13_lv_pmos
M$225 \$10 \$2 \$83 \$83 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $226 r0 *1 51.401,15.815 sg13_lv_pmos
M$226 \$64 \$95 \$220 \$220 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $227 r0 *1 52.801,15.815 sg13_lv_pmos
M$227 \$220 \$74 \$64 \$220 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $228 r0 *1 54.201,15.815 sg13_lv_pmos
M$228 \$74 \$64 \$220 \$220 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $229 r0 *1 55.601,15.815 sg13_lv_pmos
M$229 \$220 \$95 \$74 \$220 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $230 r0 *1 59.122,6.196 sg13_lv_pmos
M$230 \$48 \$9 \$49 \$220 sg13_lv_pmos W=5.999999999999998 L=0.12999999999999998
* device instance $233 r0 *1 58.259,15.815 sg13_lv_pmos
M$233 \$67 \$74 \$83 \$83 sg13_lv_pmos W=3.999999999999999 L=0.12999999999999998
* device instance $234 r0 *1 59.659,15.815 sg13_lv_pmos
M$234 \$83 \$68 \$67 \$83 sg13_lv_pmos W=3.999999999999999 L=0.12999999999999998
* device instance $235 r0 *1 61.059,15.815 sg13_lv_pmos
M$235 \$68 \$67 \$83 \$83 sg13_lv_pmos W=3.999999999999999 L=0.12999999999999998
* device instance $236 r0 *1 62.459,15.815 sg13_lv_pmos
M$236 \$83 \$64 \$68 \$83 sg13_lv_pmos W=3.999999999999999 L=0.12999999999999998
* device instance $237 r0 *1 1.445,20.146 sg13_lv_pmos
M$237 \$83 \$137 \$96 \$83 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $239 r0 *1 2.935,33.986 sg13_lv_pmos
M$239 \$187 \$36 \$83 \$83 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $240 r0 *1 3.475,34.126 sg13_lv_pmos
M$240 \$83 \$95 \$188 \$83 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $241 r0 *1 3.985,34.126 sg13_lv_pmos
M$241 \$188 \$187 \$83 \$83 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $242 r0 *1 3.365,20.146 sg13_lv_pmos
M$242 \$83 \$96 \$138 \$83 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $244 r0 *1 5.35,20.146 sg13_lv_pmos
M$244 \$83 \$92 \$140 \$83 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $246 r0 *1 6.38,20.146 sg13_lv_pmos
M$246 \$83 \$138 \$140 \$83 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $248 r0 *1 8.155,20.146 sg13_lv_pmos
M$248 \$83 \$140 \$141 \$83 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $252 r0 *1 11.035,20.146 sg13_lv_pmos
M$252 \$83 \$141 \$142 \$83 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $256 r0 *1 13.915,20.146 sg13_lv_pmos
M$256 \$83 \$142 \$143 \$83 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $260 r0 *1 16.795,20.146 sg13_lv_pmos
M$260 \$83 \$143 \$144 \$83 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $264 r0 *1 19.675,20.146 sg13_lv_pmos
M$264 \$83 \$144 \$145 \$83 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $268 r0 *1 22.555,20.146 sg13_lv_pmos
M$268 \$83 \$145 \$146 \$83 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $272 r0 *1 25.51,20.146 sg13_lv_pmos
M$272 \$83 \$146 \$148 \$83 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $274 r0 *1 26.54,20.146 sg13_lv_pmos
M$274 \$83 \$144 \$148 \$83 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $276 r0 *1 28.315,20.146 sg13_lv_pmos
M$276 \$83 \$148 \$149 \$83 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $280 r0 *1 31.135,20.146 sg13_lv_pmos
M$280 \$83 \$149 \$150 \$83 sg13_lv_pmos W=8.959999999999999
+ L=0.12999999999999995
* device instance $288 r0 *1 37.935,33.986 sg13_lv_pmos
M$288 \$193 \$19 \$83 \$83 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $289 r0 *1 38.475,34.126 sg13_lv_pmos
M$289 \$83 \$150 \$194 \$83 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $290 r0 *1 38.985,34.126 sg13_lv_pmos
M$290 \$194 \$193 \$83 \$83 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $291 r0 *1 1.51,34.141 sg13_lv_pmos
M$291 \$83 \$150 \$186 \$83 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $292 r0 *1 5.785,34.266 sg13_lv_pmos
M$292 \$83 \$95 \$189 \$83 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $293 r0 *1 6.295,34.266 sg13_lv_pmos
M$293 \$83 \$36 \$189 \$83 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $294 r0 *1 6.805,34.126 sg13_lv_pmos
M$294 \$83 \$189 \$190 \$83 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $295 r0 *1 22.577,36.411 sg13_lv_pmos
M$295 \$197 \$212 \$220 \$220 sg13_lv_pmos W=10.499999999999998
+ L=1.4999999999999996
* device instance $299 r0 *1 36.51,34.141 sg13_lv_pmos
M$299 \$83 \$95 \$192 \$83 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $300 r0 *1 40.785,34.266 sg13_lv_pmos
M$300 \$83 \$150 \$195 \$83 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $301 r0 *1 41.295,34.266 sg13_lv_pmos
M$301 \$83 \$19 \$195 \$83 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $302 r0 *1 41.805,34.126 sg13_lv_pmos
M$302 \$83 \$195 \$196 \$83 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $303 r0 *1 57.577,36.411 sg13_lv_pmos
M$303 \$48 \$213 \$220 \$220 sg13_lv_pmos W=10.499999999999998
+ L=1.4999999999999996
* device instance $307 r0 *1 10.927,36.426 sg13_lv_pmos
M$307 \$191 \$191 \$220 \$220 sg13_lv_pmos W=10.499999999999998
+ L=1.4999999999999996
* device instance $311 r0 *1 45.927,36.426 sg13_lv_pmos
M$311 \$58 \$58 \$220 \$220 sg13_lv_pmos W=10.499999999999998
+ L=1.4999999999999996
* device instance $315 r0 *1 4.41,46.621 sg13_lv_pmos
M$315 \$235 \$188 \$254 \$220 sg13_lv_pmos W=1.4999999999999998
+ L=0.12999999999999995
* device instance $316 r0 *1 6.765,46.121 sg13_lv_pmos
M$316 \$235 \$186 \$248 \$220 sg13_lv_pmos W=5.999999999999998
+ L=0.12999999999999998
* device instance $319 r0 *1 39.41,46.621 sg13_lv_pmos
M$319 \$249 \$194 \$254 \$220 sg13_lv_pmos W=1.4999999999999998
+ L=0.12999999999999995
* device instance $320 r0 *1 41.765,46.121 sg13_lv_pmos
M$320 \$249 \$192 \$197 \$220 sg13_lv_pmos W=5.999999999999998
+ L=0.12999999999999998
* device instance $323 r0 *1 43.164,9.38 cap_cmim
C$323 \$49 sub! cap_cmim w=5.77 l=5.77 m=1
* device instance $324 r0 *1 0.955,37.616 cap_cmim
C$324 \$236 \$235 cap_cmim w=5.77 l=5.77 m=1
* device instance $325 r0 *1 35.955,37.616 cap_cmim
C$325 \$246 \$249 cap_cmim w=5.77 l=5.77 m=1
* device instance $326 r0 *1 9.56,39.436 cap_cmim
C$326 \$212 \$236 cap_cmim w=8.16 l=8.16 m=1
* device instance $327 r0 *1 44.56,39.436 cap_cmim
C$327 \$213 \$246 cap_cmim w=8.16 l=8.16 m=1
* device instance $328 r0 *1 20.88,39.441 cap_cmim
C$328 \$197 \$247 cap_cmim w=8.16 l=8.16 m=1
* device instance $329 r0 *1 55.88,39.441 cap_cmim
C$329 \$48 \$237 cap_cmim w=8.16 l=8.16 m=1
.ENDS IDSM2_T4

* Extracted by KLayout with SG13G2 LVS runset on : 06/05/2024 00:42

* cell integ_5_split2.1
* pin sub!
.SUBCKT integ_5_split2.1 sub!
* device instance $1 r0 *1 3.05,0.289 sg13_lv_nmos
M$1 \$4 \$11 \$3 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $2 r0 *1 -4.112,0.291 sg13_lv_pmos
M$2 \$3 \$1 \$4 \$2 sg13_lv_pmos W=6.0 L=0.12999999999999998
.ENDS integ_5_split2.1

* Extracted by KLayout with SG13G2 LVS runset on : 03/05/2024 04:45

* cell sg13g2_Clamp_P8N8D
.SUBCKT sg13g2_Clamp_P8N8D
* device instance $1 r0 *1 34.58,6.08 sg13_hv_pmos
M$1 \$3 \$11 \$6 \$3 sg13_hv_pmos W=26.639999999999993 L=0.5999999999999999
* device instance $3 r0 *1 37.6,6.08 sg13_hv_pmos
M$3 \$3 \$11 \$7 \$3 sg13_hv_pmos W=26.639999999999993 L=0.5999999999999999
* device instance $5 r0 *1 40.62,6.08 sg13_hv_pmos
M$5 \$3 \$11 \$8 \$3 sg13_hv_pmos W=26.639999999999993 L=0.5999999999999999
* device instance $7 r0 *1 43.64,6.08 sg13_hv_pmos
M$7 \$3 \$11 \$9 \$3 sg13_hv_pmos W=26.639999999999993 L=0.5999999999999999
* device instance $17 r0 *1 17.975,16.19 dpantenna
D$17 \$11 \$3 dpantenna A=0.192 P=1.88 m=1
.ENDS sg13g2_Clamp_P8N8D

* Extracted by KLayout with SG13G2 LVS runset on : 03/05/2024 04:42

* cell sg13g2_GateLevelUpInv
* pin sub!
.SUBCKT sg13g2_GateLevelUpInv sub!
* device instance $1 r0 *1 0.51,-8.995 sg13_lv_nmos
M$1 \$12 \$11 sub! sub! sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $2 r0 *1 4.02,-8.995 sg13_lv_nmos
M$2 \$13 \$11 sub! sub! sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $3 r0 *1 0.67,-12.68 sg13_hv_nmos
M$3 \$5 \$11 sub! sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $4 r0 *1 1.5,-12.68 sg13_hv_nmos
M$4 sub! \$12 \$6 sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $5 r0 *1 2.84,-12.68 sg13_hv_nmos
M$5 sub! \$6 \$2 sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $6 r0 *1 4.18,-12.68 sg13_hv_nmos
M$6 \$7 \$11 sub! sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $7 r0 *1 5.01,-12.68 sg13_hv_nmos
M$7 sub! \$13 \$8 sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $8 r0 *1 6.35,-12.68 sg13_hv_nmos
M$8 sub! \$8 \$3 sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $9 r0 *1 0.51,-4.005 sg13_lv_pmos
M$9 \$12 \$11 \$26 \$26 sg13_lv_pmos W=4.749999999999999 L=0.12999999999999998
* device instance $10 r0 *1 4.02,-4.005 sg13_lv_pmos
M$10 \$13 \$11 \$26 \$26 sg13_lv_pmos W=4.749999999999999 L=0.12999999999999998
* device instance $11 r0 *1 0.67,-16.82 sg13_hv_pmos
M$11 \$5 \$6 \$1 \$1 sg13_hv_pmos W=0.29999999999999993 L=0.44999999999999984
* device instance $12 r0 *1 1.5,-16.82 sg13_hv_pmos
M$12 \$1 \$5 \$6 \$1 sg13_hv_pmos W=0.29999999999999993 L=0.44999999999999984
* device instance $13 r0 *1 4.18,-16.82 sg13_hv_pmos
M$13 \$7 \$8 \$1 \$1 sg13_hv_pmos W=0.29999999999999993 L=0.44999999999999984
* device instance $14 r0 *1 5.01,-16.82 sg13_hv_pmos
M$14 \$1 \$7 \$8 \$1 sg13_hv_pmos W=0.29999999999999993 L=0.44999999999999984
* device instance $15 r0 *1 2.84,-16.82 sg13_hv_pmos
M$15 \$1 \$6 \$2 \$1 sg13_hv_pmos W=3.899999999999999 L=0.4499999999999999
* device instance $16 r0 *1 6.35,-16.82 sg13_hv_pmos
M$16 \$1 \$8 \$3 \$1 sg13_hv_pmos W=3.899999999999999 L=0.4499999999999999
.ENDS sg13g2_GateLevelUpInv

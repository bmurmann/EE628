* Extracted by KLayout with SG13G2 LVS runset on : 09/05/2024 14:31

* cell comp_5_splitTop
* pin Q_N
* pin Q
* pin VDD
* pin D
* pin sub!
.SUBCKT comp_5_splitTop Q_N Q VDD D sub!
* device instance $1 r0 *1 -5.365,-1.685 sg13_lv_nmos
M$1 \$16 D \$31 sub! sg13_lv_nmos W=0.42 L=0.13
* device instance $2 r0 *1 -5.055,-1.685 sg13_lv_nmos
M$2 \$31 \$8 sub! sub! sg13_lv_nmos W=0.42 L=0.13
* device instance $3 r0 *1 -4.475,-1.3 sg13_lv_nmos
M$3 sub! \$39 \$9 sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $4 r0 *1 3.365,-1.685 sg13_lv_nmos
M$4 \$18 \$20 sub! sub! sg13_lv_nmos W=0.42 L=0.13
* device instance $5 r0 *1 3.875,-1.685 sg13_lv_nmos
M$5 sub! \$8 \$36 sub! sg13_lv_nmos W=0.42 L=0.13
* device instance $6 r0 *1 4.185,-1.685 sg13_lv_nmos
M$6 \$36 \$19 \$20 sub! sg13_lv_nmos W=0.42 L=0.13
* device instance $7 r0 *1 -3.385,-1.62 sg13_lv_nmos
M$7 sub! \$8 \$33 sub! sg13_lv_nmos W=0.42 L=0.13
* device instance $8 r0 *1 -3.075,-1.62 sg13_lv_nmos
M$8 \$33 \$9 \$17 sub! sg13_lv_nmos W=0.42 L=0.13
* device instance $9 r0 *1 22.37,-2.276 sg13_lv_nmos
M$9 sub! \$26 \$3 sub! sg13_lv_nmos W=2.0 L=1.0
* device instance $10 r0 *1 6.225,-1.575 sg13_lv_nmos
M$10 sub! \$19 \$22 sub! sg13_lv_nmos W=0.64 L=0.13
* device instance $11 r0 *1 5.205,-1.525 sg13_lv_nmos
M$11 sub! \$19 Q_N sub! sg13_lv_nmos W=1.48 L=0.13
* device instance $13 r0 *1 7.245,-1.525 sg13_lv_nmos
M$13 sub! \$22 Q sub! sg13_lv_nmos W=1.48 L=0.13
* device instance $15 r0 *1 -8.365,-1.505 sg13_lv_nmos
M$15 sub! \$38 \$15 sub! sg13_lv_nmos W=1.48 L=0.13
* device instance $17 r0 *1 -7.345,-1.455 sg13_lv_nmos
M$17 sub! D \$38 sub! sg13_lv_nmos W=0.64 L=0.13
* device instance $18 r0 *1 10.016,-1.505 sg13_lv_nmos
M$18 sub! \$40 \$8 sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $19 r0 *1 11.451,-1.505 sg13_lv_nmos
M$19 sub! \$4 \$24 sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $20 r0 *1 1.78,-1.3 sg13_lv_nmos
M$20 \$19 \$10 \$18 sub! sg13_lv_nmos W=0.42 L=0.13
* device instance $21 r0 *1 2.315,-1.46 sg13_lv_nmos
M$21 \$9 \$53 \$19 sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $22 r0 *1 -0.53,-1.42 sg13_lv_nmos
M$22 sub! \$10 \$53 sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $23 r0 *1 0.57,-1.42 sg13_lv_nmos
M$23 sub! \$4 \$10 sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $24 r0 *1 -2.3,-0.895 sg13_lv_nmos
M$24 \$16 \$10 \$39 sub! sg13_lv_nmos W=0.42 L=0.13
* device instance $25 r0 *1 -1.79,-0.895 sg13_lv_nmos
M$25 \$39 \$53 \$17 sub! sg13_lv_nmos W=0.42 L=0.13
* device instance $26 r0 *1 25.73,-0.609 sg13_lv_nmos
M$26 \$5 \$54 \$27 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $27 r0 *1 27.375,-0.609 sg13_lv_nmos
M$27 \$27 \$55 \$3 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $28 r0 *1 -7.497,2.424 sg13_lv_nmos
M$28 sub! \$54 \$79 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $29 r0 *1 12.004,3.106 sg13_lv_nmos
M$29 \$26 \$4 \$25 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $30 r0 *1 22.37,3.385 sg13_lv_nmos
M$30 sub! \$95 \$64 sub! sg13_lv_nmos W=2.0 L=1.0
* device instance $31 r0 *1 25.73,5.052 sg13_lv_nmos
M$31 \$54 \$5 \$83 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $32 r0 *1 27.375,5.052 sg13_lv_nmos
M$32 \$83 \$55 \$64 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $33 r0 *1 -7.455,5.923 sg13_lv_nmos
M$33 D \$113 \$79 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $34 r0 *1 -7.497,8.224 sg13_lv_nmos
M$34 sub! \$5 \$100 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $35 r0 *1 -7.455,11.723 sg13_lv_nmos
M$35 \$113 D \$100 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $36 r0 *1 2.725,-0.11 sg13_lv_pmos
M$36 \$19 \$53 \$61 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $37 r0 *1 3.105,-0.11 sg13_lv_pmos
M$37 \$61 \$20 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $38 r0 *1 3.715,-0.11 sg13_lv_pmos
M$38 VDD \$8 \$20 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $39 r0 *1 4.225,-0.11 sg13_lv_pmos
M$39 VDD \$19 \$20 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $40 r0 *1 5.785,-0.005 sg13_lv_pmos
M$40 VDD \$19 \$22 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $41 r0 *1 4.765,0.055 sg13_lv_pmos
M$41 VDD \$19 Q_N VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $43 r0 *1 2.03,0.18 sg13_lv_pmos
M$43 \$9 \$10 \$19 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $44 r0 *1 -5.475,-0.095 sg13_lv_pmos
M$44 VDD D \$16 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $45 r0 *1 -4.965,-0.095 sg13_lv_pmos
M$45 VDD \$8 \$16 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $46 r0 *1 -4.515,0.195 sg13_lv_pmos
M$46 VDD \$39 \$9 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $47 r0 *1 23.879,-1.583 sg13_lv_pmos
M$47 \$2 \$54 \$5 \$2 sg13_lv_pmos W=4.0 L=0.13
* device instance $48 r0 *1 29.226,-1.583 sg13_lv_pmos
M$48 \$5 \$55 \$2 \$2 sg13_lv_pmos W=4.0 L=0.13
* device instance $49 r0 *1 -3.465,0.27 sg13_lv_pmos
M$49 \$39 \$8 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $50 r0 *1 -2.73,0.27 sg13_lv_pmos
M$50 VDD \$9 \$58 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $51 r0 *1 -2.34,0.27 sg13_lv_pmos
M$51 \$58 \$10 \$39 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $52 r0 *1 -1.83,0.27 sg13_lv_pmos
M$52 \$39 \$53 \$16 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $53 r0 *1 -0.13,0.145 sg13_lv_pmos
M$53 \$53 \$10 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $54 r0 *1 0.595,0.145 sg13_lv_pmos
M$54 VDD \$4 \$10 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $55 r0 *1 -7.345,0.17 sg13_lv_pmos
M$55 VDD D \$38 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $56 r0 *1 -8.365,0.155 sg13_lv_pmos
M$56 VDD \$38 \$15 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $58 r0 *1 6.87,0.155 sg13_lv_pmos
M$58 VDD \$22 Q VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $60 r0 *1 10.026,0.17 sg13_lv_pmos
M$60 VDD \$40 \$8 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $61 r0 *1 11.461,0.17 sg13_lv_pmos
M$61 VDD \$4 \$24 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $62 r0 *1 13.289,1.106 sg13_lv_pmos
M$62 \$25 \$24 \$26 \$2 sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $63 r0 *1 23.879,4.078 sg13_lv_pmos
M$63 \$2 \$5 \$54 \$2 sg13_lv_pmos W=4.0 L=0.13
* device instance $64 r0 *1 29.226,4.078 sg13_lv_pmos
M$64 \$54 \$55 \$2 \$2 sg13_lv_pmos W=4.0 L=0.13
* device instance $65 r0 *1 -8.755,5.288 sg13_lv_pmos
M$65 D \$54 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $66 r0 *1 -5.313,5.288 sg13_lv_pmos
M$66 VDD \$113 D VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $67 r0 *1 -8.755,11.088 sg13_lv_pmos
M$67 \$113 \$5 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $68 r0 *1 -5.313,11.088 sg13_lv_pmos
M$68 VDD D \$113 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $69 r0 *1 13.778,-2.645 cap_cmim
C$69 \$26 sub! cap_cmim w=5.77 l=5.77 m=1
.ENDS comp_5_splitTop

* Extracted by KLayout with SG13G2 LVS runset on : 01/05/2024 23:06

* cell padring
.SUBCKT padring
* device instance $1 r0 *1 240.255,159.005 sg13_lv_nmos
M$1 res_c \$186 IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $2 r0 *1 440.255,159.005 sg13_lv_nmos
M$2 ck4_c \$187 IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $3 r0 *1 540.255,159.005 sg13_lv_nmos
M$3 ck5_c \$188 IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $4 r0 *1 640.255,159.005 sg13_lv_nmos
M$4 ck6_c \$189 IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $5 r0 *1 800.995,217.48 sg13_lv_nmos
M$5 \$237 out6_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $6 r0 *1 800.995,220.99 sg13_lv_nmos
M$6 \$264 out6_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $7 r0 *1 800.995,317.48 sg13_lv_nmos
M$7 \$350 out5_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $8 r0 *1 800.995,320.99 sg13_lv_nmos
M$8 \$377 out5_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $9 r0 *1 800.995,417.48 sg13_lv_nmos
M$9 \$463 out4_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $10 r0 *1 800.995,420.99 sg13_lv_nmos
M$10 \$490 out4_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $11 r0 *1 800.995,717.48 sg13_lv_nmos
M$11 \$750 out3_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $12 r0 *1 800.995,720.99 sg13_lv_nmos
M$12 \$777 out3_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $13 r0 *1 800.995,817.48 sg13_lv_nmos
M$13 \$863 out2_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $14 r0 *1 800.995,820.99 sg13_lv_nmos
M$14 \$890 out2_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $15 r0 *1 800.995,917.48 sg13_lv_nmos
M$15 \$976 out1_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $16 r0 *1 800.995,920.99 sg13_lv_nmos
M$16 \$1003 out1_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $17 r0 *1 440.255,980.995 sg13_lv_nmos
M$17 ck3_c \$1067 IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $18 r0 *1 540.255,980.995 sg13_lv_nmos
M$18 ck2_c \$1068 IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $19 r0 *1 640.255,980.995 sg13_lv_nmos
M$19 ck1_c \$1069 IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $20 r0 *1 241.765,159.055 sg13_hv_nmos
M$20 IOVSS|VSS \$129 \$186 IOVSS|VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $21 r0 *1 441.765,159.055 sg13_hv_nmos
M$21 IOVSS|VSS \$130 \$187 IOVSS|VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $22 r0 *1 541.765,159.055 sg13_hv_nmos
M$22 IOVSS|VSS \$132 \$188 IOVSS|VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $23 r0 *1 641.765,159.055 sg13_hv_nmos
M$23 IOVSS|VSS \$133 \$189 IOVSS|VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $24 r0 *1 -169.05,205.52 sg13_hv_nmos
M$24 IOVSS|VSS \$227 IN6|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $25 r0 *1 -169.05,207.3 sg13_hv_nmos
M$25 IN6|PAD \$227 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $26 r0 *1 -169.05,208.54 sg13_hv_nmos
M$26 IOVSS|VSS \$227 IN6|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $27 r0 *1 -169.05,210.32 sg13_hv_nmos
M$27 IN6|PAD \$227 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $28 r0 *1 -169.05,211.56 sg13_hv_nmos
M$28 IOVSS|VSS \$227 IN6|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $29 r0 *1 -169.05,213.34 sg13_hv_nmos
M$29 IN6|PAD \$227 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $30 r0 *1 -169.05,214.58 sg13_hv_nmos
M$30 IOVSS|VSS \$227 IN6|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $31 r0 *1 -169.05,216.36 sg13_hv_nmos
M$31 IN6|PAD \$227 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $32 r0 *1 -169.05,217.6 sg13_hv_nmos
M$32 IOVSS|VSS \$227 IN6|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $33 r0 *1 -169.05,219.38 sg13_hv_nmos
M$33 IN6|PAD \$227 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $34 r0 *1 -169.05,220.62 sg13_hv_nmos
M$34 IOVSS|VSS \$227 IN6|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $35 r0 *1 -169.05,222.4 sg13_hv_nmos
M$35 IN6|PAD \$227 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $36 r0 *1 -169.05,223.64 sg13_hv_nmos
M$36 IOVSS|VSS \$227 IN6|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $37 r0 *1 -169.05,225.42 sg13_hv_nmos
M$37 IN6|PAD \$227 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $38 r0 *1 -169.05,226.66 sg13_hv_nmos
M$38 IOVSS|VSS \$227 IN6|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $39 r0 *1 -169.05,228.44 sg13_hv_nmos
M$39 IN6|PAD \$227 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $40 r0 *1 -169.05,229.68 sg13_hv_nmos
M$40 IOVSS|VSS \$227 IN6|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $41 r0 *1 -169.05,231.46 sg13_hv_nmos
M$41 IN6|PAD \$227 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $42 r0 *1 -169.05,232.7 sg13_hv_nmos
M$42 IOVSS|VSS \$227 IN6|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $43 r0 *1 -169.05,234.48 sg13_hv_nmos
M$43 IN6|PAD \$227 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $44 r0 *1 949.05,214.58 sg13_hv_nmos
M$44 IOVSS|VSS \$253 OUT6 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $45 r0 *1 949.05,216.36 sg13_hv_nmos
M$45 OUT6 \$253 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $46 r0 *1 949.05,217.6 sg13_hv_nmos
M$46 IOVSS|VSS \$253 OUT6 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $47 r0 *1 949.05,219.38 sg13_hv_nmos
M$47 OUT6 \$253 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $48 r0 *1 949.05,220.62 sg13_hv_nmos
M$48 IOVSS|VSS \$253 OUT6 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $49 r0 *1 949.05,222.4 sg13_hv_nmos
M$49 OUT6 \$253 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $50 r0 *1 949.05,223.64 sg13_hv_nmos
M$50 IOVSS|VSS \$253 OUT6 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $51 r0 *1 949.05,225.42 sg13_hv_nmos
M$51 OUT6 \$253 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $52 r0 *1 804.68,217.64 sg13_hv_nmos
M$52 \$238 out6_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $53 r0 *1 804.68,218.47 sg13_hv_nmos
M$53 IOVSS|VSS \$237 \$248 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $54 r0 *1 804.68,219.81 sg13_hv_nmos
M$54 IOVSS|VSS \$248 \$253 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $55 r0 *1 804.68,221.15 sg13_hv_nmos
M$55 \$265 out6_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $56 r0 *1 804.68,221.98 sg13_hv_nmos
M$56 IOVSS|VSS \$264 \$272 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $57 r0 *1 804.68,223.32 sg13_hv_nmos
M$57 IOVSS|VSS \$272 \$218 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $58 r0 *1 -169.05,305.52 sg13_hv_nmos
M$58 IOVSS|VSS \$340 IN5|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $59 r0 *1 -169.05,307.3 sg13_hv_nmos
M$59 IN5|PAD \$340 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $60 r0 *1 -169.05,308.54 sg13_hv_nmos
M$60 IOVSS|VSS \$340 IN5|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $61 r0 *1 -169.05,310.32 sg13_hv_nmos
M$61 IN5|PAD \$340 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $62 r0 *1 -169.05,311.56 sg13_hv_nmos
M$62 IOVSS|VSS \$340 IN5|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $63 r0 *1 -169.05,313.34 sg13_hv_nmos
M$63 IN5|PAD \$340 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $64 r0 *1 -169.05,314.58 sg13_hv_nmos
M$64 IOVSS|VSS \$340 IN5|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $65 r0 *1 -169.05,316.36 sg13_hv_nmos
M$65 IN5|PAD \$340 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $66 r0 *1 -169.05,317.6 sg13_hv_nmos
M$66 IOVSS|VSS \$340 IN5|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $67 r0 *1 -169.05,319.38 sg13_hv_nmos
M$67 IN5|PAD \$340 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $68 r0 *1 -169.05,320.62 sg13_hv_nmos
M$68 IOVSS|VSS \$340 IN5|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $69 r0 *1 -169.05,322.4 sg13_hv_nmos
M$69 IN5|PAD \$340 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $70 r0 *1 -169.05,323.64 sg13_hv_nmos
M$70 IOVSS|VSS \$340 IN5|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $71 r0 *1 -169.05,325.42 sg13_hv_nmos
M$71 IN5|PAD \$340 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $72 r0 *1 -169.05,326.66 sg13_hv_nmos
M$72 IOVSS|VSS \$340 IN5|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $73 r0 *1 -169.05,328.44 sg13_hv_nmos
M$73 IN5|PAD \$340 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $74 r0 *1 -169.05,329.68 sg13_hv_nmos
M$74 IOVSS|VSS \$340 IN5|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $75 r0 *1 -169.05,331.46 sg13_hv_nmos
M$75 IN5|PAD \$340 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $76 r0 *1 -169.05,332.7 sg13_hv_nmos
M$76 IOVSS|VSS \$340 IN5|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $77 r0 *1 -169.05,334.48 sg13_hv_nmos
M$77 IN5|PAD \$340 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $78 r0 *1 949.05,314.58 sg13_hv_nmos
M$78 IOVSS|VSS \$366 OUT5 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $79 r0 *1 949.05,316.36 sg13_hv_nmos
M$79 OUT5 \$366 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $80 r0 *1 949.05,317.6 sg13_hv_nmos
M$80 IOVSS|VSS \$366 OUT5 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $81 r0 *1 949.05,319.38 sg13_hv_nmos
M$81 OUT5 \$366 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $82 r0 *1 949.05,320.62 sg13_hv_nmos
M$82 IOVSS|VSS \$366 OUT5 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $83 r0 *1 949.05,322.4 sg13_hv_nmos
M$83 OUT5 \$366 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $84 r0 *1 949.05,323.64 sg13_hv_nmos
M$84 IOVSS|VSS \$366 OUT5 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $85 r0 *1 949.05,325.42 sg13_hv_nmos
M$85 OUT5 \$366 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $86 r0 *1 804.68,317.64 sg13_hv_nmos
M$86 \$351 out5_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $87 r0 *1 804.68,318.47 sg13_hv_nmos
M$87 IOVSS|VSS \$350 \$361 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $88 r0 *1 804.68,319.81 sg13_hv_nmos
M$88 IOVSS|VSS \$361 \$366 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $89 r0 *1 804.68,321.15 sg13_hv_nmos
M$89 \$378 out5_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $90 r0 *1 804.68,321.98 sg13_hv_nmos
M$90 IOVSS|VSS \$377 \$385 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $91 r0 *1 804.68,323.32 sg13_hv_nmos
M$91 IOVSS|VSS \$385 \$331 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $92 r0 *1 -169.05,405.52 sg13_hv_nmos
M$92 IOVSS|VSS \$453 IN4|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $93 r0 *1 -169.05,407.3 sg13_hv_nmos
M$93 IN4|PAD \$453 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $94 r0 *1 -169.05,408.54 sg13_hv_nmos
M$94 IOVSS|VSS \$453 IN4|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $95 r0 *1 -169.05,410.32 sg13_hv_nmos
M$95 IN4|PAD \$453 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $96 r0 *1 -169.05,411.56 sg13_hv_nmos
M$96 IOVSS|VSS \$453 IN4|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $97 r0 *1 -169.05,413.34 sg13_hv_nmos
M$97 IN4|PAD \$453 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $98 r0 *1 -169.05,414.58 sg13_hv_nmos
M$98 IOVSS|VSS \$453 IN4|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $99 r0 *1 -169.05,416.36 sg13_hv_nmos
M$99 IN4|PAD \$453 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $100 r0 *1 -169.05,417.6 sg13_hv_nmos
M$100 IOVSS|VSS \$453 IN4|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $101 r0 *1 -169.05,419.38 sg13_hv_nmos
M$101 IN4|PAD \$453 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $102 r0 *1 -169.05,420.62 sg13_hv_nmos
M$102 IOVSS|VSS \$453 IN4|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $103 r0 *1 -169.05,422.4 sg13_hv_nmos
M$103 IN4|PAD \$453 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $104 r0 *1 -169.05,423.64 sg13_hv_nmos
M$104 IOVSS|VSS \$453 IN4|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $105 r0 *1 -169.05,425.42 sg13_hv_nmos
M$105 IN4|PAD \$453 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $106 r0 *1 -169.05,426.66 sg13_hv_nmos
M$106 IOVSS|VSS \$453 IN4|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $107 r0 *1 -169.05,428.44 sg13_hv_nmos
M$107 IN4|PAD \$453 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $108 r0 *1 -169.05,429.68 sg13_hv_nmos
M$108 IOVSS|VSS \$453 IN4|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $109 r0 *1 -169.05,431.46 sg13_hv_nmos
M$109 IN4|PAD \$453 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $110 r0 *1 -169.05,432.7 sg13_hv_nmos
M$110 IOVSS|VSS \$453 IN4|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $111 r0 *1 -169.05,434.48 sg13_hv_nmos
M$111 IN4|PAD \$453 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $112 r0 *1 949.05,414.58 sg13_hv_nmos
M$112 IOVSS|VSS \$479 OUT4 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $113 r0 *1 949.05,416.36 sg13_hv_nmos
M$113 OUT4 \$479 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $114 r0 *1 949.05,417.6 sg13_hv_nmos
M$114 IOVSS|VSS \$479 OUT4 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $115 r0 *1 949.05,419.38 sg13_hv_nmos
M$115 OUT4 \$479 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $116 r0 *1 949.05,420.62 sg13_hv_nmos
M$116 IOVSS|VSS \$479 OUT4 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $117 r0 *1 949.05,422.4 sg13_hv_nmos
M$117 OUT4 \$479 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $118 r0 *1 949.05,423.64 sg13_hv_nmos
M$118 IOVSS|VSS \$479 OUT4 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $119 r0 *1 949.05,425.42 sg13_hv_nmos
M$119 OUT4 \$479 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $120 r0 *1 804.68,417.64 sg13_hv_nmos
M$120 \$464 out4_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $121 r0 *1 804.68,418.47 sg13_hv_nmos
M$121 IOVSS|VSS \$463 \$474 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $122 r0 *1 804.68,419.81 sg13_hv_nmos
M$122 IOVSS|VSS \$474 \$479 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $123 r0 *1 804.68,421.15 sg13_hv_nmos
M$123 \$491 out4_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $124 r0 *1 804.68,421.98 sg13_hv_nmos
M$124 IOVSS|VSS \$490 \$498 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $125 r0 *1 804.68,423.32 sg13_hv_nmos
M$125 IOVSS|VSS \$498 \$444 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $126 r0 *1 -169.05,505.52 sg13_hv_nmos
M$126 IOVSS|VSS \$568 PAD|VLO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $127 r0 *1 -169.05,507.3 sg13_hv_nmos
M$127 PAD|VLO \$568 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $128 r0 *1 -169.05,508.54 sg13_hv_nmos
M$128 IOVSS|VSS \$568 PAD|VLO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $129 r0 *1 -169.05,510.32 sg13_hv_nmos
M$129 PAD|VLO \$568 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $130 r0 *1 -169.05,511.56 sg13_hv_nmos
M$130 IOVSS|VSS \$568 PAD|VLO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $131 r0 *1 -169.05,513.34 sg13_hv_nmos
M$131 PAD|VLO \$568 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $132 r0 *1 -169.05,514.58 sg13_hv_nmos
M$132 IOVSS|VSS \$568 PAD|VLO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $133 r0 *1 -169.05,516.36 sg13_hv_nmos
M$133 PAD|VLO \$568 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $134 r0 *1 -169.05,517.6 sg13_hv_nmos
M$134 IOVSS|VSS \$568 PAD|VLO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $135 r0 *1 -169.05,519.38 sg13_hv_nmos
M$135 PAD|VLO \$568 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $136 r0 *1 -169.05,520.62 sg13_hv_nmos
M$136 IOVSS|VSS \$568 PAD|VLO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $137 r0 *1 -169.05,522.4 sg13_hv_nmos
M$137 PAD|VLO \$568 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $138 r0 *1 -169.05,523.64 sg13_hv_nmos
M$138 IOVSS|VSS \$568 PAD|VLO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $139 r0 *1 -169.05,525.42 sg13_hv_nmos
M$139 PAD|VLO \$568 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $140 r0 *1 -169.05,526.66 sg13_hv_nmos
M$140 IOVSS|VSS \$568 PAD|VLO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $141 r0 *1 -169.05,528.44 sg13_hv_nmos
M$141 PAD|VLO \$568 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $142 r0 *1 -169.05,529.68 sg13_hv_nmos
M$142 IOVSS|VSS \$568 PAD|VLO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $143 r0 *1 -169.05,531.46 sg13_hv_nmos
M$143 PAD|VLO \$568 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $144 r0 *1 -169.05,532.7 sg13_hv_nmos
M$144 IOVSS|VSS \$568 PAD|VLO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $145 r0 *1 -169.05,534.48 sg13_hv_nmos
M$145 PAD|VLO \$568 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $146 r0 *1 879.21,583.22 sg13_hv_nmos
M$146 IOVSS|VSS IOVDD \$626 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $147 r0 *1 879.21,584.1 sg13_hv_nmos
M$147 \$626 IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $148 r0 *1 879.21,584.98 sg13_hv_nmos
M$148 IOVSS|VSS IOVDD \$626 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $149 r0 *1 879.21,585.86 sg13_hv_nmos
M$149 \$626 IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $150 r0 *1 879.21,586.74 sg13_hv_nmos
M$150 IOVSS|VSS IOVDD \$626 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $151 r0 *1 879.21,587.62 sg13_hv_nmos
M$151 \$626 IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $152 r0 *1 879.21,593 sg13_hv_nmos
M$152 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $153 r0 *1 879.21,602.88 sg13_hv_nmos
M$153 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $154 r0 *1 879.21,612.76 sg13_hv_nmos
M$154 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $155 r0 *1 879.21,622.64 sg13_hv_nmos
M$155 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $156 r0 *1 879.21,632.52 sg13_hv_nmos
M$156 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $157 r0 *1 879.21,642.4 sg13_hv_nmos
M$157 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $158 r0 *1 879.21,652.28 sg13_hv_nmos
M$158 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $159 r0 *1 888.46,583.22 sg13_hv_nmos
M$159 IOVSS|VSS IOVDD \$626 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $160 r0 *1 888.46,584.1 sg13_hv_nmos
M$160 \$626 IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $161 r0 *1 888.46,584.98 sg13_hv_nmos
M$161 IOVSS|VSS IOVDD \$626 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $162 r0 *1 888.46,585.86 sg13_hv_nmos
M$162 \$626 IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $163 r0 *1 888.46,586.74 sg13_hv_nmos
M$163 IOVSS|VSS IOVDD \$626 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $164 r0 *1 888.46,587.62 sg13_hv_nmos
M$164 \$626 IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $165 r0 *1 888.46,593 sg13_hv_nmos
M$165 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $166 r0 *1 888.46,602.88 sg13_hv_nmos
M$166 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $167 r0 *1 888.46,612.76 sg13_hv_nmos
M$167 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $168 r0 *1 888.46,622.64 sg13_hv_nmos
M$168 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $169 r0 *1 888.46,632.52 sg13_hv_nmos
M$169 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $170 r0 *1 888.46,642.4 sg13_hv_nmos
M$170 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $171 r0 *1 888.46,652.28 sg13_hv_nmos
M$171 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $172 r0 *1 934.53,588.155 sg13_hv_nmos
M$172 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $173 r0 *1 934.53,589.935 sg13_hv_nmos
M$173 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $174 r0 *1 934.53,591.175 sg13_hv_nmos
M$174 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $175 r0 *1 934.53,592.955 sg13_hv_nmos
M$175 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $176 r0 *1 934.53,594.195 sg13_hv_nmos
M$176 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $177 r0 *1 934.53,595.975 sg13_hv_nmos
M$177 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $178 r0 *1 934.53,597.215 sg13_hv_nmos
M$178 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $179 r0 *1 934.53,598.995 sg13_hv_nmos
M$179 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $180 r0 *1 934.53,600.235 sg13_hv_nmos
M$180 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $181 r0 *1 934.53,602.015 sg13_hv_nmos
M$181 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $182 r0 *1 934.53,603.255 sg13_hv_nmos
M$182 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $183 r0 *1 934.53,605.035 sg13_hv_nmos
M$183 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $184 r0 *1 934.53,606.275 sg13_hv_nmos
M$184 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $185 r0 *1 934.53,608.055 sg13_hv_nmos
M$185 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $186 r0 *1 934.53,609.295 sg13_hv_nmos
M$186 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $187 r0 *1 934.53,611.075 sg13_hv_nmos
M$187 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $188 r0 *1 934.53,612.315 sg13_hv_nmos
M$188 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $189 r0 *1 934.53,614.095 sg13_hv_nmos
M$189 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $190 r0 *1 934.53,615.335 sg13_hv_nmos
M$190 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $191 r0 *1 934.53,617.115 sg13_hv_nmos
M$191 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $192 r0 *1 934.53,618.355 sg13_hv_nmos
M$192 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $193 r0 *1 934.53,620.135 sg13_hv_nmos
M$193 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $194 r0 *1 934.53,621.375 sg13_hv_nmos
M$194 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $195 r0 *1 934.53,623.155 sg13_hv_nmos
M$195 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $196 r0 *1 934.53,624.395 sg13_hv_nmos
M$196 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $197 r0 *1 934.53,626.175 sg13_hv_nmos
M$197 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $198 r0 *1 934.53,627.415 sg13_hv_nmos
M$198 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $199 r0 *1 934.53,629.195 sg13_hv_nmos
M$199 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $200 r0 *1 934.53,630.435 sg13_hv_nmos
M$200 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $201 r0 *1 934.53,632.215 sg13_hv_nmos
M$201 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $202 r0 *1 934.53,633.455 sg13_hv_nmos
M$202 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $203 r0 *1 934.53,635.235 sg13_hv_nmos
M$203 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $204 r0 *1 934.53,636.475 sg13_hv_nmos
M$204 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $205 r0 *1 934.53,638.255 sg13_hv_nmos
M$205 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $206 r0 *1 934.53,639.495 sg13_hv_nmos
M$206 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $207 r0 *1 934.53,641.275 sg13_hv_nmos
M$207 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $208 r0 *1 934.53,642.515 sg13_hv_nmos
M$208 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $209 r0 *1 934.53,644.295 sg13_hv_nmos
M$209 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $210 r0 *1 934.53,645.535 sg13_hv_nmos
M$210 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $211 r0 *1 934.53,647.315 sg13_hv_nmos
M$211 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $212 r0 *1 934.53,648.555 sg13_hv_nmos
M$212 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $213 r0 *1 934.53,650.335 sg13_hv_nmos
M$213 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $214 r0 *1 934.53,651.575 sg13_hv_nmos
M$214 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $215 r0 *1 939.37,588.155 sg13_hv_nmos
M$215 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $216 r0 *1 939.37,589.935 sg13_hv_nmos
M$216 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $217 r0 *1 939.37,591.175 sg13_hv_nmos
M$217 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $218 r0 *1 939.37,592.955 sg13_hv_nmos
M$218 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $219 r0 *1 939.37,594.195 sg13_hv_nmos
M$219 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $220 r0 *1 939.37,595.975 sg13_hv_nmos
M$220 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $221 r0 *1 939.37,597.215 sg13_hv_nmos
M$221 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $222 r0 *1 939.37,598.995 sg13_hv_nmos
M$222 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $223 r0 *1 939.37,600.235 sg13_hv_nmos
M$223 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $224 r0 *1 939.37,602.015 sg13_hv_nmos
M$224 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $225 r0 *1 939.37,603.255 sg13_hv_nmos
M$225 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $226 r0 *1 939.37,605.035 sg13_hv_nmos
M$226 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $227 r0 *1 939.37,606.275 sg13_hv_nmos
M$227 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $228 r0 *1 939.37,608.055 sg13_hv_nmos
M$228 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $229 r0 *1 939.37,609.295 sg13_hv_nmos
M$229 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $230 r0 *1 939.37,611.075 sg13_hv_nmos
M$230 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $231 r0 *1 939.37,612.315 sg13_hv_nmos
M$231 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $232 r0 *1 939.37,614.095 sg13_hv_nmos
M$232 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $233 r0 *1 939.37,615.335 sg13_hv_nmos
M$233 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $234 r0 *1 939.37,617.115 sg13_hv_nmos
M$234 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $235 r0 *1 939.37,618.355 sg13_hv_nmos
M$235 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $236 r0 *1 939.37,620.135 sg13_hv_nmos
M$236 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $237 r0 *1 939.37,621.375 sg13_hv_nmos
M$237 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $238 r0 *1 939.37,623.155 sg13_hv_nmos
M$238 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $239 r0 *1 939.37,624.395 sg13_hv_nmos
M$239 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $240 r0 *1 939.37,626.175 sg13_hv_nmos
M$240 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $241 r0 *1 939.37,627.415 sg13_hv_nmos
M$241 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $242 r0 *1 939.37,629.195 sg13_hv_nmos
M$242 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $243 r0 *1 939.37,630.435 sg13_hv_nmos
M$243 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $244 r0 *1 939.37,632.215 sg13_hv_nmos
M$244 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $245 r0 *1 939.37,633.455 sg13_hv_nmos
M$245 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $246 r0 *1 939.37,635.235 sg13_hv_nmos
M$246 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $247 r0 *1 939.37,636.475 sg13_hv_nmos
M$247 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $248 r0 *1 939.37,638.255 sg13_hv_nmos
M$248 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $249 r0 *1 939.37,639.495 sg13_hv_nmos
M$249 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $250 r0 *1 939.37,641.275 sg13_hv_nmos
M$250 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $251 r0 *1 939.37,642.515 sg13_hv_nmos
M$251 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $252 r0 *1 939.37,644.295 sg13_hv_nmos
M$252 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $253 r0 *1 939.37,645.535 sg13_hv_nmos
M$253 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $254 r0 *1 939.37,647.315 sg13_hv_nmos
M$254 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $255 r0 *1 939.37,648.555 sg13_hv_nmos
M$255 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $256 r0 *1 939.37,650.335 sg13_hv_nmos
M$256 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $257 r0 *1 939.37,651.575 sg13_hv_nmos
M$257 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $258 r0 *1 944.21,588.155 sg13_hv_nmos
M$258 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $259 r0 *1 944.21,589.935 sg13_hv_nmos
M$259 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $260 r0 *1 944.21,591.175 sg13_hv_nmos
M$260 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $261 r0 *1 944.21,592.955 sg13_hv_nmos
M$261 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $262 r0 *1 944.21,594.195 sg13_hv_nmos
M$262 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $263 r0 *1 944.21,595.975 sg13_hv_nmos
M$263 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $264 r0 *1 944.21,597.215 sg13_hv_nmos
M$264 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $265 r0 *1 944.21,598.995 sg13_hv_nmos
M$265 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $266 r0 *1 944.21,600.235 sg13_hv_nmos
M$266 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $267 r0 *1 944.21,602.015 sg13_hv_nmos
M$267 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $268 r0 *1 944.21,603.255 sg13_hv_nmos
M$268 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $269 r0 *1 944.21,605.035 sg13_hv_nmos
M$269 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $270 r0 *1 944.21,606.275 sg13_hv_nmos
M$270 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $271 r0 *1 944.21,608.055 sg13_hv_nmos
M$271 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $272 r0 *1 944.21,609.295 sg13_hv_nmos
M$272 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $273 r0 *1 944.21,611.075 sg13_hv_nmos
M$273 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $274 r0 *1 944.21,612.315 sg13_hv_nmos
M$274 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $275 r0 *1 944.21,614.095 sg13_hv_nmos
M$275 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $276 r0 *1 944.21,615.335 sg13_hv_nmos
M$276 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $277 r0 *1 944.21,617.115 sg13_hv_nmos
M$277 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $278 r0 *1 944.21,618.355 sg13_hv_nmos
M$278 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $279 r0 *1 944.21,620.135 sg13_hv_nmos
M$279 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $280 r0 *1 944.21,621.375 sg13_hv_nmos
M$280 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $281 r0 *1 944.21,623.155 sg13_hv_nmos
M$281 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $282 r0 *1 944.21,624.395 sg13_hv_nmos
M$282 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $283 r0 *1 944.21,626.175 sg13_hv_nmos
M$283 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $284 r0 *1 944.21,627.415 sg13_hv_nmos
M$284 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $285 r0 *1 944.21,629.195 sg13_hv_nmos
M$285 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $286 r0 *1 944.21,630.435 sg13_hv_nmos
M$286 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $287 r0 *1 944.21,632.215 sg13_hv_nmos
M$287 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $288 r0 *1 944.21,633.455 sg13_hv_nmos
M$288 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $289 r0 *1 944.21,635.235 sg13_hv_nmos
M$289 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $290 r0 *1 944.21,636.475 sg13_hv_nmos
M$290 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $291 r0 *1 944.21,638.255 sg13_hv_nmos
M$291 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $292 r0 *1 944.21,639.495 sg13_hv_nmos
M$292 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $293 r0 *1 944.21,641.275 sg13_hv_nmos
M$293 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $294 r0 *1 944.21,642.515 sg13_hv_nmos
M$294 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $295 r0 *1 944.21,644.295 sg13_hv_nmos
M$295 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $296 r0 *1 944.21,645.535 sg13_hv_nmos
M$296 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $297 r0 *1 944.21,647.315 sg13_hv_nmos
M$297 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $298 r0 *1 944.21,648.555 sg13_hv_nmos
M$298 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $299 r0 *1 944.21,650.335 sg13_hv_nmos
M$299 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $300 r0 *1 944.21,651.575 sg13_hv_nmos
M$300 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $301 r0 *1 949.05,588.155 sg13_hv_nmos
M$301 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $302 r0 *1 949.05,589.935 sg13_hv_nmos
M$302 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $303 r0 *1 949.05,591.175 sg13_hv_nmos
M$303 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $304 r0 *1 949.05,592.955 sg13_hv_nmos
M$304 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $305 r0 *1 949.05,594.195 sg13_hv_nmos
M$305 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $306 r0 *1 949.05,595.975 sg13_hv_nmos
M$306 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $307 r0 *1 949.05,597.215 sg13_hv_nmos
M$307 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $308 r0 *1 949.05,598.995 sg13_hv_nmos
M$308 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $309 r0 *1 949.05,600.235 sg13_hv_nmos
M$309 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $310 r0 *1 949.05,602.015 sg13_hv_nmos
M$310 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $311 r0 *1 949.05,603.255 sg13_hv_nmos
M$311 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $312 r0 *1 949.05,605.035 sg13_hv_nmos
M$312 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $313 r0 *1 949.05,606.275 sg13_hv_nmos
M$313 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $314 r0 *1 949.05,608.055 sg13_hv_nmos
M$314 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $315 r0 *1 949.05,609.295 sg13_hv_nmos
M$315 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $316 r0 *1 949.05,611.075 sg13_hv_nmos
M$316 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $317 r0 *1 949.05,612.315 sg13_hv_nmos
M$317 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $318 r0 *1 949.05,614.095 sg13_hv_nmos
M$318 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $319 r0 *1 949.05,615.335 sg13_hv_nmos
M$319 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $320 r0 *1 949.05,617.115 sg13_hv_nmos
M$320 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $321 r0 *1 949.05,618.355 sg13_hv_nmos
M$321 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $322 r0 *1 949.05,620.135 sg13_hv_nmos
M$322 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $323 r0 *1 949.05,621.375 sg13_hv_nmos
M$323 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $324 r0 *1 949.05,623.155 sg13_hv_nmos
M$324 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $325 r0 *1 949.05,624.395 sg13_hv_nmos
M$325 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $326 r0 *1 949.05,626.175 sg13_hv_nmos
M$326 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $327 r0 *1 949.05,627.415 sg13_hv_nmos
M$327 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $328 r0 *1 949.05,629.195 sg13_hv_nmos
M$328 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $329 r0 *1 949.05,630.435 sg13_hv_nmos
M$329 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $330 r0 *1 949.05,632.215 sg13_hv_nmos
M$330 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $331 r0 *1 949.05,633.455 sg13_hv_nmos
M$331 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $332 r0 *1 949.05,635.235 sg13_hv_nmos
M$332 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $333 r0 *1 949.05,636.475 sg13_hv_nmos
M$333 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $334 r0 *1 949.05,638.255 sg13_hv_nmos
M$334 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $335 r0 *1 949.05,639.495 sg13_hv_nmos
M$335 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $336 r0 *1 949.05,641.275 sg13_hv_nmos
M$336 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $337 r0 *1 949.05,642.515 sg13_hv_nmos
M$337 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $338 r0 *1 949.05,644.295 sg13_hv_nmos
M$338 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $339 r0 *1 949.05,645.535 sg13_hv_nmos
M$339 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $340 r0 *1 949.05,647.315 sg13_hv_nmos
M$340 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $341 r0 *1 949.05,648.555 sg13_hv_nmos
M$341 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $342 r0 *1 949.05,650.335 sg13_hv_nmos
M$342 IOVDD \$626 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $343 r0 *1 949.05,651.575 sg13_hv_nmos
M$343 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $344 r0 *1 -169.05,605.52 sg13_hv_nmos
M$344 IOVSS|VSS \$638 PAD|VHI IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $345 r0 *1 -169.05,607.3 sg13_hv_nmos
M$345 PAD|VHI \$638 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $346 r0 *1 -169.05,608.54 sg13_hv_nmos
M$346 IOVSS|VSS \$638 PAD|VHI IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $347 r0 *1 -169.05,610.32 sg13_hv_nmos
M$347 PAD|VHI \$638 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $348 r0 *1 -169.05,611.56 sg13_hv_nmos
M$348 IOVSS|VSS \$638 PAD|VHI IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $349 r0 *1 -169.05,613.34 sg13_hv_nmos
M$349 PAD|VHI \$638 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $350 r0 *1 -169.05,614.58 sg13_hv_nmos
M$350 IOVSS|VSS \$638 PAD|VHI IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $351 r0 *1 -169.05,616.36 sg13_hv_nmos
M$351 PAD|VHI \$638 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $352 r0 *1 -169.05,617.6 sg13_hv_nmos
M$352 IOVSS|VSS \$638 PAD|VHI IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $353 r0 *1 -169.05,619.38 sg13_hv_nmos
M$353 PAD|VHI \$638 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $354 r0 *1 -169.05,620.62 sg13_hv_nmos
M$354 IOVSS|VSS \$638 PAD|VHI IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $355 r0 *1 -169.05,622.4 sg13_hv_nmos
M$355 PAD|VHI \$638 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $356 r0 *1 -169.05,623.64 sg13_hv_nmos
M$356 IOVSS|VSS \$638 PAD|VHI IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $357 r0 *1 -169.05,625.42 sg13_hv_nmos
M$357 PAD|VHI \$638 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $358 r0 *1 -169.05,626.66 sg13_hv_nmos
M$358 IOVSS|VSS \$638 PAD|VHI IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $359 r0 *1 -169.05,628.44 sg13_hv_nmos
M$359 PAD|VHI \$638 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $360 r0 *1 -169.05,629.68 sg13_hv_nmos
M$360 IOVSS|VSS \$638 PAD|VHI IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $361 r0 *1 -169.05,631.46 sg13_hv_nmos
M$361 PAD|VHI \$638 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $362 r0 *1 -169.05,632.7 sg13_hv_nmos
M$362 IOVSS|VSS \$638 PAD|VHI IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $363 r0 *1 -169.05,634.48 sg13_hv_nmos
M$363 PAD|VHI \$638 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $364 r0 *1 -169.05,705.52 sg13_hv_nmos
M$364 IOVSS|VSS \$740 IN3|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $365 r0 *1 -169.05,707.3 sg13_hv_nmos
M$365 IN3|PAD \$740 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $366 r0 *1 -169.05,708.54 sg13_hv_nmos
M$366 IOVSS|VSS \$740 IN3|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $367 r0 *1 -169.05,710.32 sg13_hv_nmos
M$367 IN3|PAD \$740 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $368 r0 *1 -169.05,711.56 sg13_hv_nmos
M$368 IOVSS|VSS \$740 IN3|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $369 r0 *1 -169.05,713.34 sg13_hv_nmos
M$369 IN3|PAD \$740 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $370 r0 *1 -169.05,714.58 sg13_hv_nmos
M$370 IOVSS|VSS \$740 IN3|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $371 r0 *1 -169.05,716.36 sg13_hv_nmos
M$371 IN3|PAD \$740 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $372 r0 *1 -169.05,717.6 sg13_hv_nmos
M$372 IOVSS|VSS \$740 IN3|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $373 r0 *1 -169.05,719.38 sg13_hv_nmos
M$373 IN3|PAD \$740 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $374 r0 *1 -169.05,720.62 sg13_hv_nmos
M$374 IOVSS|VSS \$740 IN3|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $375 r0 *1 -169.05,722.4 sg13_hv_nmos
M$375 IN3|PAD \$740 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $376 r0 *1 -169.05,723.64 sg13_hv_nmos
M$376 IOVSS|VSS \$740 IN3|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $377 r0 *1 -169.05,725.42 sg13_hv_nmos
M$377 IN3|PAD \$740 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $378 r0 *1 -169.05,726.66 sg13_hv_nmos
M$378 IOVSS|VSS \$740 IN3|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $379 r0 *1 -169.05,728.44 sg13_hv_nmos
M$379 IN3|PAD \$740 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $380 r0 *1 -169.05,729.68 sg13_hv_nmos
M$380 IOVSS|VSS \$740 IN3|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $381 r0 *1 -169.05,731.46 sg13_hv_nmos
M$381 IN3|PAD \$740 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $382 r0 *1 -169.05,732.7 sg13_hv_nmos
M$382 IOVSS|VSS \$740 IN3|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $383 r0 *1 -169.05,734.48 sg13_hv_nmos
M$383 IN3|PAD \$740 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $384 r0 *1 949.05,714.58 sg13_hv_nmos
M$384 IOVSS|VSS \$766 OUT3 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $385 r0 *1 949.05,716.36 sg13_hv_nmos
M$385 OUT3 \$766 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $386 r0 *1 949.05,717.6 sg13_hv_nmos
M$386 IOVSS|VSS \$766 OUT3 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $387 r0 *1 949.05,719.38 sg13_hv_nmos
M$387 OUT3 \$766 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $388 r0 *1 949.05,720.62 sg13_hv_nmos
M$388 IOVSS|VSS \$766 OUT3 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $389 r0 *1 949.05,722.4 sg13_hv_nmos
M$389 OUT3 \$766 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $390 r0 *1 949.05,723.64 sg13_hv_nmos
M$390 IOVSS|VSS \$766 OUT3 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $391 r0 *1 949.05,725.42 sg13_hv_nmos
M$391 OUT3 \$766 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $392 r0 *1 804.68,717.64 sg13_hv_nmos
M$392 \$751 out3_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $393 r0 *1 804.68,718.47 sg13_hv_nmos
M$393 IOVSS|VSS \$750 \$761 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $394 r0 *1 804.68,719.81 sg13_hv_nmos
M$394 IOVSS|VSS \$761 \$766 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $395 r0 *1 804.68,721.15 sg13_hv_nmos
M$395 \$778 out3_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $396 r0 *1 804.68,721.98 sg13_hv_nmos
M$396 IOVSS|VSS \$777 \$785 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $397 r0 *1 804.68,723.32 sg13_hv_nmos
M$397 IOVSS|VSS \$785 \$731 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $398 r0 *1 -169.05,805.52 sg13_hv_nmos
M$398 IOVSS|VSS \$853 IN2|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $399 r0 *1 -169.05,807.3 sg13_hv_nmos
M$399 IN2|PAD \$853 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $400 r0 *1 -169.05,808.54 sg13_hv_nmos
M$400 IOVSS|VSS \$853 IN2|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $401 r0 *1 -169.05,810.32 sg13_hv_nmos
M$401 IN2|PAD \$853 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $402 r0 *1 -169.05,811.56 sg13_hv_nmos
M$402 IOVSS|VSS \$853 IN2|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $403 r0 *1 -169.05,813.34 sg13_hv_nmos
M$403 IN2|PAD \$853 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $404 r0 *1 -169.05,814.58 sg13_hv_nmos
M$404 IOVSS|VSS \$853 IN2|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $405 r0 *1 -169.05,816.36 sg13_hv_nmos
M$405 IN2|PAD \$853 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $406 r0 *1 -169.05,817.6 sg13_hv_nmos
M$406 IOVSS|VSS \$853 IN2|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $407 r0 *1 -169.05,819.38 sg13_hv_nmos
M$407 IN2|PAD \$853 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $408 r0 *1 -169.05,820.62 sg13_hv_nmos
M$408 IOVSS|VSS \$853 IN2|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $409 r0 *1 -169.05,822.4 sg13_hv_nmos
M$409 IN2|PAD \$853 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $410 r0 *1 -169.05,823.64 sg13_hv_nmos
M$410 IOVSS|VSS \$853 IN2|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $411 r0 *1 -169.05,825.42 sg13_hv_nmos
M$411 IN2|PAD \$853 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $412 r0 *1 -169.05,826.66 sg13_hv_nmos
M$412 IOVSS|VSS \$853 IN2|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $413 r0 *1 -169.05,828.44 sg13_hv_nmos
M$413 IN2|PAD \$853 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $414 r0 *1 -169.05,829.68 sg13_hv_nmos
M$414 IOVSS|VSS \$853 IN2|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $415 r0 *1 -169.05,831.46 sg13_hv_nmos
M$415 IN2|PAD \$853 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $416 r0 *1 -169.05,832.7 sg13_hv_nmos
M$416 IOVSS|VSS \$853 IN2|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $417 r0 *1 -169.05,834.48 sg13_hv_nmos
M$417 IN2|PAD \$853 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $418 r0 *1 949.05,814.58 sg13_hv_nmos
M$418 IOVSS|VSS \$879 OUT2 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $419 r0 *1 949.05,816.36 sg13_hv_nmos
M$419 OUT2 \$879 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $420 r0 *1 949.05,817.6 sg13_hv_nmos
M$420 IOVSS|VSS \$879 OUT2 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $421 r0 *1 949.05,819.38 sg13_hv_nmos
M$421 OUT2 \$879 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $422 r0 *1 949.05,820.62 sg13_hv_nmos
M$422 IOVSS|VSS \$879 OUT2 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $423 r0 *1 949.05,822.4 sg13_hv_nmos
M$423 OUT2 \$879 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $424 r0 *1 949.05,823.64 sg13_hv_nmos
M$424 IOVSS|VSS \$879 OUT2 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $425 r0 *1 949.05,825.42 sg13_hv_nmos
M$425 OUT2 \$879 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $426 r0 *1 804.68,817.64 sg13_hv_nmos
M$426 \$864 out2_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $427 r0 *1 804.68,818.47 sg13_hv_nmos
M$427 IOVSS|VSS \$863 \$874 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $428 r0 *1 804.68,819.81 sg13_hv_nmos
M$428 IOVSS|VSS \$874 \$879 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $429 r0 *1 804.68,821.15 sg13_hv_nmos
M$429 \$891 out2_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $430 r0 *1 804.68,821.98 sg13_hv_nmos
M$430 IOVSS|VSS \$890 \$898 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $431 r0 *1 804.68,823.32 sg13_hv_nmos
M$431 IOVSS|VSS \$898 \$844 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $432 r0 *1 -169.05,905.52 sg13_hv_nmos
M$432 IOVSS|VSS \$966 IN1|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $433 r0 *1 -169.05,907.3 sg13_hv_nmos
M$433 IN1|PAD \$966 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $434 r0 *1 -169.05,908.54 sg13_hv_nmos
M$434 IOVSS|VSS \$966 IN1|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $435 r0 *1 -169.05,910.32 sg13_hv_nmos
M$435 IN1|PAD \$966 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $436 r0 *1 -169.05,911.56 sg13_hv_nmos
M$436 IOVSS|VSS \$966 IN1|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $437 r0 *1 -169.05,913.34 sg13_hv_nmos
M$437 IN1|PAD \$966 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $438 r0 *1 -169.05,914.58 sg13_hv_nmos
M$438 IOVSS|VSS \$966 IN1|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $439 r0 *1 -169.05,916.36 sg13_hv_nmos
M$439 IN1|PAD \$966 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $440 r0 *1 -169.05,917.6 sg13_hv_nmos
M$440 IOVSS|VSS \$966 IN1|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $441 r0 *1 -169.05,919.38 sg13_hv_nmos
M$441 IN1|PAD \$966 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $442 r0 *1 -169.05,920.62 sg13_hv_nmos
M$442 IOVSS|VSS \$966 IN1|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $443 r0 *1 -169.05,922.4 sg13_hv_nmos
M$443 IN1|PAD \$966 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $444 r0 *1 -169.05,923.64 sg13_hv_nmos
M$444 IOVSS|VSS \$966 IN1|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $445 r0 *1 -169.05,925.42 sg13_hv_nmos
M$445 IN1|PAD \$966 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $446 r0 *1 -169.05,926.66 sg13_hv_nmos
M$446 IOVSS|VSS \$966 IN1|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $447 r0 *1 -169.05,928.44 sg13_hv_nmos
M$447 IN1|PAD \$966 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $448 r0 *1 -169.05,929.68 sg13_hv_nmos
M$448 IOVSS|VSS \$966 IN1|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $449 r0 *1 -169.05,931.46 sg13_hv_nmos
M$449 IN1|PAD \$966 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $450 r0 *1 -169.05,932.7 sg13_hv_nmos
M$450 IOVSS|VSS \$966 IN1|PAD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $451 r0 *1 -169.05,934.48 sg13_hv_nmos
M$451 IN1|PAD \$966 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $452 r0 *1 949.05,914.58 sg13_hv_nmos
M$452 IOVSS|VSS \$992 OUT1 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $453 r0 *1 949.05,916.36 sg13_hv_nmos
M$453 OUT1 \$992 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $454 r0 *1 949.05,917.6 sg13_hv_nmos
M$454 IOVSS|VSS \$992 OUT1 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $455 r0 *1 949.05,919.38 sg13_hv_nmos
M$455 OUT1 \$992 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $456 r0 *1 949.05,920.62 sg13_hv_nmos
M$456 IOVSS|VSS \$992 OUT1 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $457 r0 *1 949.05,922.4 sg13_hv_nmos
M$457 OUT1 \$992 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $458 r0 *1 949.05,923.64 sg13_hv_nmos
M$458 IOVSS|VSS \$992 OUT1 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $459 r0 *1 949.05,925.42 sg13_hv_nmos
M$459 OUT1 \$992 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $460 r0 *1 804.68,917.64 sg13_hv_nmos
M$460 \$977 out1_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $461 r0 *1 804.68,918.47 sg13_hv_nmos
M$461 IOVSS|VSS \$976 \$987 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $462 r0 *1 804.68,919.81 sg13_hv_nmos
M$462 IOVSS|VSS \$987 \$992 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $463 r0 *1 804.68,921.15 sg13_hv_nmos
M$463 \$1004 out1_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $464 r0 *1 804.68,921.98 sg13_hv_nmos
M$464 IOVSS|VSS \$1003 \$1011 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $465 r0 *1 804.68,923.32 sg13_hv_nmos
M$465 IOVSS|VSS \$1011 \$957 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $466 r0 *1 441.765,980.945 sg13_hv_nmos
M$466 IOVSS|VSS \$1070 \$1067 IOVSS|VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $467 r0 *1 541.765,980.945 sg13_hv_nmos
M$467 IOVSS|VSS \$1071 \$1068 IOVSS|VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $468 r0 *1 641.765,980.945 sg13_hv_nmos
M$468 IOVSS|VSS \$1072 \$1069 IOVSS|VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $469 r0 *1 3.22,1059.21 sg13_hv_nmos
M$469 IOVSS|VSS AVDD|IOVDD \$1143 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $470 r0 *1 4.1,1059.21 sg13_hv_nmos
M$470 \$1143 AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $471 r0 *1 4.98,1059.21 sg13_hv_nmos
M$471 IOVSS|VSS AVDD|IOVDD \$1143 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $472 r0 *1 5.86,1059.21 sg13_hv_nmos
M$472 \$1143 AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $473 r0 *1 6.74,1059.21 sg13_hv_nmos
M$473 IOVSS|VSS AVDD|IOVDD \$1143 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $474 r0 *1 7.62,1059.21 sg13_hv_nmos
M$474 \$1143 AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $475 r0 *1 13,1059.21 sg13_hv_nmos
M$475 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $476 r0 *1 22.88,1059.21 sg13_hv_nmos
M$476 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $477 r0 *1 32.76,1059.21 sg13_hv_nmos
M$477 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $478 r0 *1 42.64,1059.21 sg13_hv_nmos
M$478 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $479 r0 *1 52.52,1059.21 sg13_hv_nmos
M$479 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $480 r0 *1 62.4,1059.21 sg13_hv_nmos
M$480 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $481 r0 *1 72.28,1059.21 sg13_hv_nmos
M$481 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $482 r0 *1 303.22,1059.21 sg13_hv_nmos
M$482 IOVSS|VSS IOVDD \$1144 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $483 r0 *1 304.1,1059.21 sg13_hv_nmos
M$483 \$1144 IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $484 r0 *1 304.98,1059.21 sg13_hv_nmos
M$484 IOVSS|VSS IOVDD \$1144 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $485 r0 *1 305.86,1059.21 sg13_hv_nmos
M$485 \$1144 IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $486 r0 *1 306.74,1059.21 sg13_hv_nmos
M$486 IOVSS|VSS IOVDD \$1144 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $487 r0 *1 307.62,1059.21 sg13_hv_nmos
M$487 \$1144 IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $488 r0 *1 313,1059.21 sg13_hv_nmos
M$488 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $489 r0 *1 322.88,1059.21 sg13_hv_nmos
M$489 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $490 r0 *1 332.76,1059.21 sg13_hv_nmos
M$490 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $491 r0 *1 342.64,1059.21 sg13_hv_nmos
M$491 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $492 r0 *1 352.52,1059.21 sg13_hv_nmos
M$492 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $493 r0 *1 362.4,1059.21 sg13_hv_nmos
M$493 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $494 r0 *1 372.28,1059.21 sg13_hv_nmos
M$494 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $495 r0 *1 703.22,1059.21 sg13_hv_nmos
M$495 IOVSS|VSS VDD \$1145 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $496 r0 *1 704.1,1059.21 sg13_hv_nmos
M$496 \$1145 VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $497 r0 *1 704.98,1059.21 sg13_hv_nmos
M$497 IOVSS|VSS VDD \$1145 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $498 r0 *1 705.86,1059.21 sg13_hv_nmos
M$498 \$1145 VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $499 r0 *1 706.74,1059.21 sg13_hv_nmos
M$499 IOVSS|VSS VDD \$1145 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $500 r0 *1 707.62,1059.21 sg13_hv_nmos
M$500 \$1145 VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $501 r0 *1 713,1059.21 sg13_hv_nmos
M$501 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $502 r0 *1 722.88,1059.21 sg13_hv_nmos
M$502 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $503 r0 *1 732.76,1059.21 sg13_hv_nmos
M$503 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $504 r0 *1 742.64,1059.21 sg13_hv_nmos
M$504 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $505 r0 *1 752.52,1059.21 sg13_hv_nmos
M$505 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $506 r0 *1 762.4,1059.21 sg13_hv_nmos
M$506 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $507 r0 *1 772.28,1059.21 sg13_hv_nmos
M$507 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $508 r0 *1 3.22,1068.46 sg13_hv_nmos
M$508 IOVSS|VSS AVDD|IOVDD \$1143 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $509 r0 *1 4.1,1068.46 sg13_hv_nmos
M$509 \$1143 AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $510 r0 *1 4.98,1068.46 sg13_hv_nmos
M$510 IOVSS|VSS AVDD|IOVDD \$1143 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $511 r0 *1 5.86,1068.46 sg13_hv_nmos
M$511 \$1143 AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $512 r0 *1 6.74,1068.46 sg13_hv_nmos
M$512 IOVSS|VSS AVDD|IOVDD \$1143 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $513 r0 *1 7.62,1068.46 sg13_hv_nmos
M$513 \$1143 AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $514 r0 *1 13,1068.46 sg13_hv_nmos
M$514 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $515 r0 *1 22.88,1068.46 sg13_hv_nmos
M$515 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $516 r0 *1 32.76,1068.46 sg13_hv_nmos
M$516 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $517 r0 *1 42.64,1068.46 sg13_hv_nmos
M$517 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $518 r0 *1 52.52,1068.46 sg13_hv_nmos
M$518 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $519 r0 *1 62.4,1068.46 sg13_hv_nmos
M$519 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $520 r0 *1 72.28,1068.46 sg13_hv_nmos
M$520 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $521 r0 *1 303.22,1068.46 sg13_hv_nmos
M$521 IOVSS|VSS IOVDD \$1144 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $522 r0 *1 304.1,1068.46 sg13_hv_nmos
M$522 \$1144 IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $523 r0 *1 304.98,1068.46 sg13_hv_nmos
M$523 IOVSS|VSS IOVDD \$1144 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $524 r0 *1 305.86,1068.46 sg13_hv_nmos
M$524 \$1144 IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $525 r0 *1 306.74,1068.46 sg13_hv_nmos
M$525 IOVSS|VSS IOVDD \$1144 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $526 r0 *1 307.62,1068.46 sg13_hv_nmos
M$526 \$1144 IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $527 r0 *1 313,1068.46 sg13_hv_nmos
M$527 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $528 r0 *1 322.88,1068.46 sg13_hv_nmos
M$528 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $529 r0 *1 332.76,1068.46 sg13_hv_nmos
M$529 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $530 r0 *1 342.64,1068.46 sg13_hv_nmos
M$530 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $531 r0 *1 352.52,1068.46 sg13_hv_nmos
M$531 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $532 r0 *1 362.4,1068.46 sg13_hv_nmos
M$532 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $533 r0 *1 372.28,1068.46 sg13_hv_nmos
M$533 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $534 r0 *1 703.22,1068.46 sg13_hv_nmos
M$534 IOVSS|VSS VDD \$1145 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $535 r0 *1 704.1,1068.46 sg13_hv_nmos
M$535 \$1145 VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $536 r0 *1 704.98,1068.46 sg13_hv_nmos
M$536 IOVSS|VSS VDD \$1145 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $537 r0 *1 705.86,1068.46 sg13_hv_nmos
M$537 \$1145 VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $538 r0 *1 706.74,1068.46 sg13_hv_nmos
M$538 IOVSS|VSS VDD \$1145 IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $539 r0 *1 707.62,1068.46 sg13_hv_nmos
M$539 \$1145 VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=0.4999999999999999
* device instance $540 r0 *1 713,1068.46 sg13_hv_nmos
M$540 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $541 r0 *1 722.88,1068.46 sg13_hv_nmos
M$541 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $542 r0 *1 732.76,1068.46 sg13_hv_nmos
M$542 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $543 r0 *1 742.64,1068.46 sg13_hv_nmos
M$543 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $544 r0 *1 752.52,1068.46 sg13_hv_nmos
M$544 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $545 r0 *1 762.4,1068.46 sg13_hv_nmos
M$545 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $546 r0 *1 772.28,1068.46 sg13_hv_nmos
M$546 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=8.999999999999998
+ L=9.499999999999996
* device instance $547 r0 *1 8.155,1114.53 sg13_hv_nmos
M$547 IOVSS|VSS \$1143 \$1316 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $548 r0 *1 9.935,1114.53 sg13_hv_nmos
M$548 \$1316 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $549 r0 *1 11.175,1114.53 sg13_hv_nmos
M$549 IOVSS|VSS \$1143 \$1317 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $550 r0 *1 12.955,1114.53 sg13_hv_nmos
M$550 \$1317 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $551 r0 *1 14.195,1114.53 sg13_hv_nmos
M$551 IOVSS|VSS \$1143 \$1318 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $552 r0 *1 15.975,1114.53 sg13_hv_nmos
M$552 \$1318 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $553 r0 *1 17.215,1114.53 sg13_hv_nmos
M$553 IOVSS|VSS \$1143 \$1319 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $554 r0 *1 18.995,1114.53 sg13_hv_nmos
M$554 \$1319 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $555 r0 *1 20.235,1114.53 sg13_hv_nmos
M$555 IOVSS|VSS \$1143 \$1320 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $556 r0 *1 22.015,1114.53 sg13_hv_nmos
M$556 \$1320 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $557 r0 *1 23.255,1114.53 sg13_hv_nmos
M$557 IOVSS|VSS \$1143 \$1321 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $558 r0 *1 25.035,1114.53 sg13_hv_nmos
M$558 \$1321 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $559 r0 *1 26.275,1114.53 sg13_hv_nmos
M$559 IOVSS|VSS \$1143 \$1322 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $560 r0 *1 28.055,1114.53 sg13_hv_nmos
M$560 \$1322 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $561 r0 *1 29.295,1114.53 sg13_hv_nmos
M$561 IOVSS|VSS \$1143 \$1323 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $562 r0 *1 31.075,1114.53 sg13_hv_nmos
M$562 \$1323 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $563 r0 *1 32.315,1114.53 sg13_hv_nmos
M$563 IOVSS|VSS \$1143 \$1324 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $564 r0 *1 34.095,1114.53 sg13_hv_nmos
M$564 \$1324 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $565 r0 *1 35.335,1114.53 sg13_hv_nmos
M$565 IOVSS|VSS \$1143 \$1325 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $566 r0 *1 37.115,1114.53 sg13_hv_nmos
M$566 \$1325 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $567 r0 *1 38.355,1114.53 sg13_hv_nmos
M$567 IOVSS|VSS \$1143 \$1326 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $568 r0 *1 40.135,1114.53 sg13_hv_nmos
M$568 \$1326 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $569 r0 *1 41.375,1114.53 sg13_hv_nmos
M$569 IOVSS|VSS \$1143 \$1327 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $570 r0 *1 43.155,1114.53 sg13_hv_nmos
M$570 \$1327 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $571 r0 *1 44.395,1114.53 sg13_hv_nmos
M$571 IOVSS|VSS \$1143 \$1328 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $572 r0 *1 46.175,1114.53 sg13_hv_nmos
M$572 \$1328 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $573 r0 *1 47.415,1114.53 sg13_hv_nmos
M$573 IOVSS|VSS \$1143 \$1329 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $574 r0 *1 49.195,1114.53 sg13_hv_nmos
M$574 \$1329 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $575 r0 *1 50.435,1114.53 sg13_hv_nmos
M$575 IOVSS|VSS \$1143 \$1330 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $576 r0 *1 52.215,1114.53 sg13_hv_nmos
M$576 \$1330 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $577 r0 *1 53.455,1114.53 sg13_hv_nmos
M$577 IOVSS|VSS \$1143 \$1331 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $578 r0 *1 55.235,1114.53 sg13_hv_nmos
M$578 \$1331 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $579 r0 *1 56.475,1114.53 sg13_hv_nmos
M$579 IOVSS|VSS \$1143 \$1332 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $580 r0 *1 58.255,1114.53 sg13_hv_nmos
M$580 \$1332 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $581 r0 *1 59.495,1114.53 sg13_hv_nmos
M$581 IOVSS|VSS \$1143 \$1333 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $582 r0 *1 61.275,1114.53 sg13_hv_nmos
M$582 \$1333 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $583 r0 *1 62.515,1114.53 sg13_hv_nmos
M$583 IOVSS|VSS \$1143 \$1334 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $584 r0 *1 64.295,1114.53 sg13_hv_nmos
M$584 \$1334 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $585 r0 *1 65.535,1114.53 sg13_hv_nmos
M$585 IOVSS|VSS \$1143 \$1335 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $586 r0 *1 67.315,1114.53 sg13_hv_nmos
M$586 \$1335 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $587 r0 *1 68.555,1114.53 sg13_hv_nmos
M$587 IOVSS|VSS \$1143 \$1336 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $588 r0 *1 70.335,1114.53 sg13_hv_nmos
M$588 \$1336 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $589 r0 *1 71.575,1114.53 sg13_hv_nmos
M$589 IOVSS|VSS \$1143 \$1337 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $590 r0 *1 308.155,1114.53 sg13_hv_nmos
M$590 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $591 r0 *1 309.935,1114.53 sg13_hv_nmos
M$591 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $592 r0 *1 311.175,1114.53 sg13_hv_nmos
M$592 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $593 r0 *1 312.955,1114.53 sg13_hv_nmos
M$593 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $594 r0 *1 314.195,1114.53 sg13_hv_nmos
M$594 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $595 r0 *1 315.975,1114.53 sg13_hv_nmos
M$595 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $596 r0 *1 317.215,1114.53 sg13_hv_nmos
M$596 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $597 r0 *1 318.995,1114.53 sg13_hv_nmos
M$597 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $598 r0 *1 320.235,1114.53 sg13_hv_nmos
M$598 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $599 r0 *1 322.015,1114.53 sg13_hv_nmos
M$599 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $600 r0 *1 323.255,1114.53 sg13_hv_nmos
M$600 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $601 r0 *1 325.035,1114.53 sg13_hv_nmos
M$601 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $602 r0 *1 326.275,1114.53 sg13_hv_nmos
M$602 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $603 r0 *1 328.055,1114.53 sg13_hv_nmos
M$603 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $604 r0 *1 329.295,1114.53 sg13_hv_nmos
M$604 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $605 r0 *1 331.075,1114.53 sg13_hv_nmos
M$605 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $606 r0 *1 332.315,1114.53 sg13_hv_nmos
M$606 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $607 r0 *1 334.095,1114.53 sg13_hv_nmos
M$607 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $608 r0 *1 335.335,1114.53 sg13_hv_nmos
M$608 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $609 r0 *1 337.115,1114.53 sg13_hv_nmos
M$609 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $610 r0 *1 338.355,1114.53 sg13_hv_nmos
M$610 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $611 r0 *1 340.135,1114.53 sg13_hv_nmos
M$611 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $612 r0 *1 341.375,1114.53 sg13_hv_nmos
M$612 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $613 r0 *1 343.155,1114.53 sg13_hv_nmos
M$613 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $614 r0 *1 344.395,1114.53 sg13_hv_nmos
M$614 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $615 r0 *1 346.175,1114.53 sg13_hv_nmos
M$615 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $616 r0 *1 347.415,1114.53 sg13_hv_nmos
M$616 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $617 r0 *1 349.195,1114.53 sg13_hv_nmos
M$617 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $618 r0 *1 350.435,1114.53 sg13_hv_nmos
M$618 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $619 r0 *1 352.215,1114.53 sg13_hv_nmos
M$619 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $620 r0 *1 353.455,1114.53 sg13_hv_nmos
M$620 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $621 r0 *1 355.235,1114.53 sg13_hv_nmos
M$621 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $622 r0 *1 356.475,1114.53 sg13_hv_nmos
M$622 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $623 r0 *1 358.255,1114.53 sg13_hv_nmos
M$623 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $624 r0 *1 359.495,1114.53 sg13_hv_nmos
M$624 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $625 r0 *1 361.275,1114.53 sg13_hv_nmos
M$625 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $626 r0 *1 362.515,1114.53 sg13_hv_nmos
M$626 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $627 r0 *1 364.295,1114.53 sg13_hv_nmos
M$627 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $628 r0 *1 365.535,1114.53 sg13_hv_nmos
M$628 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $629 r0 *1 367.315,1114.53 sg13_hv_nmos
M$629 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $630 r0 *1 368.555,1114.53 sg13_hv_nmos
M$630 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $631 r0 *1 370.335,1114.53 sg13_hv_nmos
M$631 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $632 r0 *1 371.575,1114.53 sg13_hv_nmos
M$632 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $633 r0 *1 708.155,1114.53 sg13_hv_nmos
M$633 IOVSS|VSS \$1145 \$1338 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $634 r0 *1 709.935,1114.53 sg13_hv_nmos
M$634 \$1338 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $635 r0 *1 711.175,1114.53 sg13_hv_nmos
M$635 IOVSS|VSS \$1145 \$1339 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $636 r0 *1 712.955,1114.53 sg13_hv_nmos
M$636 \$1339 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $637 r0 *1 714.195,1114.53 sg13_hv_nmos
M$637 IOVSS|VSS \$1145 \$1340 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $638 r0 *1 715.975,1114.53 sg13_hv_nmos
M$638 \$1340 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $639 r0 *1 717.215,1114.53 sg13_hv_nmos
M$639 IOVSS|VSS \$1145 \$1341 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $640 r0 *1 718.995,1114.53 sg13_hv_nmos
M$640 \$1341 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $641 r0 *1 720.235,1114.53 sg13_hv_nmos
M$641 IOVSS|VSS \$1145 \$1342 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $642 r0 *1 722.015,1114.53 sg13_hv_nmos
M$642 \$1342 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $643 r0 *1 723.255,1114.53 sg13_hv_nmos
M$643 IOVSS|VSS \$1145 \$1343 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $644 r0 *1 725.035,1114.53 sg13_hv_nmos
M$644 \$1343 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $645 r0 *1 726.275,1114.53 sg13_hv_nmos
M$645 IOVSS|VSS \$1145 \$1344 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $646 r0 *1 728.055,1114.53 sg13_hv_nmos
M$646 \$1344 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $647 r0 *1 729.295,1114.53 sg13_hv_nmos
M$647 IOVSS|VSS \$1145 \$1345 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $648 r0 *1 731.075,1114.53 sg13_hv_nmos
M$648 \$1345 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $649 r0 *1 732.315,1114.53 sg13_hv_nmos
M$649 IOVSS|VSS \$1145 \$1346 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $650 r0 *1 734.095,1114.53 sg13_hv_nmos
M$650 \$1346 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $651 r0 *1 735.335,1114.53 sg13_hv_nmos
M$651 IOVSS|VSS \$1145 \$1347 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $652 r0 *1 737.115,1114.53 sg13_hv_nmos
M$652 \$1347 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $653 r0 *1 738.355,1114.53 sg13_hv_nmos
M$653 IOVSS|VSS \$1145 \$1348 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $654 r0 *1 740.135,1114.53 sg13_hv_nmos
M$654 \$1348 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $655 r0 *1 741.375,1114.53 sg13_hv_nmos
M$655 IOVSS|VSS \$1145 \$1349 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $656 r0 *1 743.155,1114.53 sg13_hv_nmos
M$656 \$1349 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $657 r0 *1 744.395,1114.53 sg13_hv_nmos
M$657 IOVSS|VSS \$1145 \$1350 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $658 r0 *1 746.175,1114.53 sg13_hv_nmos
M$658 \$1350 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $659 r0 *1 747.415,1114.53 sg13_hv_nmos
M$659 IOVSS|VSS \$1145 \$1351 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $660 r0 *1 749.195,1114.53 sg13_hv_nmos
M$660 \$1351 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $661 r0 *1 750.435,1114.53 sg13_hv_nmos
M$661 IOVSS|VSS \$1145 \$1352 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $662 r0 *1 752.215,1114.53 sg13_hv_nmos
M$662 \$1352 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $663 r0 *1 753.455,1114.53 sg13_hv_nmos
M$663 IOVSS|VSS \$1145 \$1353 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $664 r0 *1 755.235,1114.53 sg13_hv_nmos
M$664 \$1353 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $665 r0 *1 756.475,1114.53 sg13_hv_nmos
M$665 IOVSS|VSS \$1145 \$1354 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $666 r0 *1 758.255,1114.53 sg13_hv_nmos
M$666 \$1354 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $667 r0 *1 759.495,1114.53 sg13_hv_nmos
M$667 IOVSS|VSS \$1145 \$1355 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $668 r0 *1 761.275,1114.53 sg13_hv_nmos
M$668 \$1355 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $669 r0 *1 762.515,1114.53 sg13_hv_nmos
M$669 IOVSS|VSS \$1145 \$1356 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $670 r0 *1 764.295,1114.53 sg13_hv_nmos
M$670 \$1356 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $671 r0 *1 765.535,1114.53 sg13_hv_nmos
M$671 IOVSS|VSS \$1145 \$1357 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $672 r0 *1 767.315,1114.53 sg13_hv_nmos
M$672 \$1357 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $673 r0 *1 768.555,1114.53 sg13_hv_nmos
M$673 IOVSS|VSS \$1145 \$1358 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $674 r0 *1 770.335,1114.53 sg13_hv_nmos
M$674 \$1358 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $675 r0 *1 771.575,1114.53 sg13_hv_nmos
M$675 IOVSS|VSS \$1145 \$1359 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $676 r0 *1 8.155,1119.37 sg13_hv_nmos
M$676 IOVSS|VSS \$1143 \$1316 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $677 r0 *1 9.935,1119.37 sg13_hv_nmos
M$677 \$1316 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $678 r0 *1 11.175,1119.37 sg13_hv_nmos
M$678 IOVSS|VSS \$1143 \$1317 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $679 r0 *1 12.955,1119.37 sg13_hv_nmos
M$679 \$1317 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $680 r0 *1 14.195,1119.37 sg13_hv_nmos
M$680 IOVSS|VSS \$1143 \$1318 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $681 r0 *1 15.975,1119.37 sg13_hv_nmos
M$681 \$1318 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $682 r0 *1 17.215,1119.37 sg13_hv_nmos
M$682 IOVSS|VSS \$1143 \$1319 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $683 r0 *1 18.995,1119.37 sg13_hv_nmos
M$683 \$1319 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $684 r0 *1 20.235,1119.37 sg13_hv_nmos
M$684 IOVSS|VSS \$1143 \$1320 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $685 r0 *1 22.015,1119.37 sg13_hv_nmos
M$685 \$1320 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $686 r0 *1 23.255,1119.37 sg13_hv_nmos
M$686 IOVSS|VSS \$1143 \$1321 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $687 r0 *1 25.035,1119.37 sg13_hv_nmos
M$687 \$1321 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $688 r0 *1 26.275,1119.37 sg13_hv_nmos
M$688 IOVSS|VSS \$1143 \$1322 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $689 r0 *1 28.055,1119.37 sg13_hv_nmos
M$689 \$1322 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $690 r0 *1 29.295,1119.37 sg13_hv_nmos
M$690 IOVSS|VSS \$1143 \$1323 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $691 r0 *1 31.075,1119.37 sg13_hv_nmos
M$691 \$1323 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $692 r0 *1 32.315,1119.37 sg13_hv_nmos
M$692 IOVSS|VSS \$1143 \$1324 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $693 r0 *1 34.095,1119.37 sg13_hv_nmos
M$693 \$1324 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $694 r0 *1 35.335,1119.37 sg13_hv_nmos
M$694 IOVSS|VSS \$1143 \$1325 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $695 r0 *1 37.115,1119.37 sg13_hv_nmos
M$695 \$1325 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $696 r0 *1 38.355,1119.37 sg13_hv_nmos
M$696 IOVSS|VSS \$1143 \$1326 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $697 r0 *1 40.135,1119.37 sg13_hv_nmos
M$697 \$1326 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $698 r0 *1 41.375,1119.37 sg13_hv_nmos
M$698 IOVSS|VSS \$1143 \$1327 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $699 r0 *1 43.155,1119.37 sg13_hv_nmos
M$699 \$1327 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $700 r0 *1 44.395,1119.37 sg13_hv_nmos
M$700 IOVSS|VSS \$1143 \$1328 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $701 r0 *1 46.175,1119.37 sg13_hv_nmos
M$701 \$1328 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $702 r0 *1 47.415,1119.37 sg13_hv_nmos
M$702 IOVSS|VSS \$1143 \$1329 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $703 r0 *1 49.195,1119.37 sg13_hv_nmos
M$703 \$1329 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $704 r0 *1 50.435,1119.37 sg13_hv_nmos
M$704 IOVSS|VSS \$1143 \$1330 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $705 r0 *1 52.215,1119.37 sg13_hv_nmos
M$705 \$1330 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $706 r0 *1 53.455,1119.37 sg13_hv_nmos
M$706 IOVSS|VSS \$1143 \$1331 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $707 r0 *1 55.235,1119.37 sg13_hv_nmos
M$707 \$1331 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $708 r0 *1 56.475,1119.37 sg13_hv_nmos
M$708 IOVSS|VSS \$1143 \$1332 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $709 r0 *1 58.255,1119.37 sg13_hv_nmos
M$709 \$1332 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $710 r0 *1 59.495,1119.37 sg13_hv_nmos
M$710 IOVSS|VSS \$1143 \$1333 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $711 r0 *1 61.275,1119.37 sg13_hv_nmos
M$711 \$1333 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $712 r0 *1 62.515,1119.37 sg13_hv_nmos
M$712 IOVSS|VSS \$1143 \$1334 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $713 r0 *1 64.295,1119.37 sg13_hv_nmos
M$713 \$1334 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $714 r0 *1 65.535,1119.37 sg13_hv_nmos
M$714 IOVSS|VSS \$1143 \$1335 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $715 r0 *1 67.315,1119.37 sg13_hv_nmos
M$715 \$1335 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $716 r0 *1 68.555,1119.37 sg13_hv_nmos
M$716 IOVSS|VSS \$1143 \$1336 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $717 r0 *1 70.335,1119.37 sg13_hv_nmos
M$717 \$1336 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $718 r0 *1 71.575,1119.37 sg13_hv_nmos
M$718 IOVSS|VSS \$1143 \$1337 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $719 r0 *1 308.155,1119.37 sg13_hv_nmos
M$719 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $720 r0 *1 309.935,1119.37 sg13_hv_nmos
M$720 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $721 r0 *1 311.175,1119.37 sg13_hv_nmos
M$721 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $722 r0 *1 312.955,1119.37 sg13_hv_nmos
M$722 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $723 r0 *1 314.195,1119.37 sg13_hv_nmos
M$723 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $724 r0 *1 315.975,1119.37 sg13_hv_nmos
M$724 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $725 r0 *1 317.215,1119.37 sg13_hv_nmos
M$725 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $726 r0 *1 318.995,1119.37 sg13_hv_nmos
M$726 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $727 r0 *1 320.235,1119.37 sg13_hv_nmos
M$727 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $728 r0 *1 322.015,1119.37 sg13_hv_nmos
M$728 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $729 r0 *1 323.255,1119.37 sg13_hv_nmos
M$729 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $730 r0 *1 325.035,1119.37 sg13_hv_nmos
M$730 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $731 r0 *1 326.275,1119.37 sg13_hv_nmos
M$731 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $732 r0 *1 328.055,1119.37 sg13_hv_nmos
M$732 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $733 r0 *1 329.295,1119.37 sg13_hv_nmos
M$733 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $734 r0 *1 331.075,1119.37 sg13_hv_nmos
M$734 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $735 r0 *1 332.315,1119.37 sg13_hv_nmos
M$735 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $736 r0 *1 334.095,1119.37 sg13_hv_nmos
M$736 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $737 r0 *1 335.335,1119.37 sg13_hv_nmos
M$737 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $738 r0 *1 337.115,1119.37 sg13_hv_nmos
M$738 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $739 r0 *1 338.355,1119.37 sg13_hv_nmos
M$739 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $740 r0 *1 340.135,1119.37 sg13_hv_nmos
M$740 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $741 r0 *1 341.375,1119.37 sg13_hv_nmos
M$741 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $742 r0 *1 343.155,1119.37 sg13_hv_nmos
M$742 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $743 r0 *1 344.395,1119.37 sg13_hv_nmos
M$743 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $744 r0 *1 346.175,1119.37 sg13_hv_nmos
M$744 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $745 r0 *1 347.415,1119.37 sg13_hv_nmos
M$745 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $746 r0 *1 349.195,1119.37 sg13_hv_nmos
M$746 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $747 r0 *1 350.435,1119.37 sg13_hv_nmos
M$747 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $748 r0 *1 352.215,1119.37 sg13_hv_nmos
M$748 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $749 r0 *1 353.455,1119.37 sg13_hv_nmos
M$749 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $750 r0 *1 355.235,1119.37 sg13_hv_nmos
M$750 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $751 r0 *1 356.475,1119.37 sg13_hv_nmos
M$751 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $752 r0 *1 358.255,1119.37 sg13_hv_nmos
M$752 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $753 r0 *1 359.495,1119.37 sg13_hv_nmos
M$753 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $754 r0 *1 361.275,1119.37 sg13_hv_nmos
M$754 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $755 r0 *1 362.515,1119.37 sg13_hv_nmos
M$755 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $756 r0 *1 364.295,1119.37 sg13_hv_nmos
M$756 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $757 r0 *1 365.535,1119.37 sg13_hv_nmos
M$757 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $758 r0 *1 367.315,1119.37 sg13_hv_nmos
M$758 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $759 r0 *1 368.555,1119.37 sg13_hv_nmos
M$759 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $760 r0 *1 370.335,1119.37 sg13_hv_nmos
M$760 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $761 r0 *1 371.575,1119.37 sg13_hv_nmos
M$761 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $762 r0 *1 708.155,1119.37 sg13_hv_nmos
M$762 IOVSS|VSS \$1145 \$1338 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $763 r0 *1 709.935,1119.37 sg13_hv_nmos
M$763 \$1338 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $764 r0 *1 711.175,1119.37 sg13_hv_nmos
M$764 IOVSS|VSS \$1145 \$1339 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $765 r0 *1 712.955,1119.37 sg13_hv_nmos
M$765 \$1339 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $766 r0 *1 714.195,1119.37 sg13_hv_nmos
M$766 IOVSS|VSS \$1145 \$1340 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $767 r0 *1 715.975,1119.37 sg13_hv_nmos
M$767 \$1340 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $768 r0 *1 717.215,1119.37 sg13_hv_nmos
M$768 IOVSS|VSS \$1145 \$1341 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $769 r0 *1 718.995,1119.37 sg13_hv_nmos
M$769 \$1341 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $770 r0 *1 720.235,1119.37 sg13_hv_nmos
M$770 IOVSS|VSS \$1145 \$1342 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $771 r0 *1 722.015,1119.37 sg13_hv_nmos
M$771 \$1342 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $772 r0 *1 723.255,1119.37 sg13_hv_nmos
M$772 IOVSS|VSS \$1145 \$1343 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $773 r0 *1 725.035,1119.37 sg13_hv_nmos
M$773 \$1343 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $774 r0 *1 726.275,1119.37 sg13_hv_nmos
M$774 IOVSS|VSS \$1145 \$1344 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $775 r0 *1 728.055,1119.37 sg13_hv_nmos
M$775 \$1344 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $776 r0 *1 729.295,1119.37 sg13_hv_nmos
M$776 IOVSS|VSS \$1145 \$1345 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $777 r0 *1 731.075,1119.37 sg13_hv_nmos
M$777 \$1345 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $778 r0 *1 732.315,1119.37 sg13_hv_nmos
M$778 IOVSS|VSS \$1145 \$1346 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $779 r0 *1 734.095,1119.37 sg13_hv_nmos
M$779 \$1346 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $780 r0 *1 735.335,1119.37 sg13_hv_nmos
M$780 IOVSS|VSS \$1145 \$1347 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $781 r0 *1 737.115,1119.37 sg13_hv_nmos
M$781 \$1347 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $782 r0 *1 738.355,1119.37 sg13_hv_nmos
M$782 IOVSS|VSS \$1145 \$1348 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $783 r0 *1 740.135,1119.37 sg13_hv_nmos
M$783 \$1348 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $784 r0 *1 741.375,1119.37 sg13_hv_nmos
M$784 IOVSS|VSS \$1145 \$1349 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $785 r0 *1 743.155,1119.37 sg13_hv_nmos
M$785 \$1349 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $786 r0 *1 744.395,1119.37 sg13_hv_nmos
M$786 IOVSS|VSS \$1145 \$1350 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $787 r0 *1 746.175,1119.37 sg13_hv_nmos
M$787 \$1350 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $788 r0 *1 747.415,1119.37 sg13_hv_nmos
M$788 IOVSS|VSS \$1145 \$1351 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $789 r0 *1 749.195,1119.37 sg13_hv_nmos
M$789 \$1351 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $790 r0 *1 750.435,1119.37 sg13_hv_nmos
M$790 IOVSS|VSS \$1145 \$1352 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $791 r0 *1 752.215,1119.37 sg13_hv_nmos
M$791 \$1352 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $792 r0 *1 753.455,1119.37 sg13_hv_nmos
M$792 IOVSS|VSS \$1145 \$1353 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $793 r0 *1 755.235,1119.37 sg13_hv_nmos
M$793 \$1353 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $794 r0 *1 756.475,1119.37 sg13_hv_nmos
M$794 IOVSS|VSS \$1145 \$1354 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $795 r0 *1 758.255,1119.37 sg13_hv_nmos
M$795 \$1354 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $796 r0 *1 759.495,1119.37 sg13_hv_nmos
M$796 IOVSS|VSS \$1145 \$1355 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $797 r0 *1 761.275,1119.37 sg13_hv_nmos
M$797 \$1355 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $798 r0 *1 762.515,1119.37 sg13_hv_nmos
M$798 IOVSS|VSS \$1145 \$1356 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $799 r0 *1 764.295,1119.37 sg13_hv_nmos
M$799 \$1356 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $800 r0 *1 765.535,1119.37 sg13_hv_nmos
M$800 IOVSS|VSS \$1145 \$1357 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $801 r0 *1 767.315,1119.37 sg13_hv_nmos
M$801 \$1357 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $802 r0 *1 768.555,1119.37 sg13_hv_nmos
M$802 IOVSS|VSS \$1145 \$1358 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $803 r0 *1 770.335,1119.37 sg13_hv_nmos
M$803 \$1358 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $804 r0 *1 771.575,1119.37 sg13_hv_nmos
M$804 IOVSS|VSS \$1145 \$1359 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $805 r0 *1 8.155,1124.21 sg13_hv_nmos
M$805 IOVSS|VSS \$1143 \$1316 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $806 r0 *1 9.935,1124.21 sg13_hv_nmos
M$806 \$1316 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $807 r0 *1 11.175,1124.21 sg13_hv_nmos
M$807 IOVSS|VSS \$1143 \$1317 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $808 r0 *1 12.955,1124.21 sg13_hv_nmos
M$808 \$1317 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $809 r0 *1 14.195,1124.21 sg13_hv_nmos
M$809 IOVSS|VSS \$1143 \$1318 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $810 r0 *1 15.975,1124.21 sg13_hv_nmos
M$810 \$1318 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $811 r0 *1 17.215,1124.21 sg13_hv_nmos
M$811 IOVSS|VSS \$1143 \$1319 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $812 r0 *1 18.995,1124.21 sg13_hv_nmos
M$812 \$1319 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $813 r0 *1 20.235,1124.21 sg13_hv_nmos
M$813 IOVSS|VSS \$1143 \$1320 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $814 r0 *1 22.015,1124.21 sg13_hv_nmos
M$814 \$1320 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $815 r0 *1 23.255,1124.21 sg13_hv_nmos
M$815 IOVSS|VSS \$1143 \$1321 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $816 r0 *1 25.035,1124.21 sg13_hv_nmos
M$816 \$1321 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $817 r0 *1 26.275,1124.21 sg13_hv_nmos
M$817 IOVSS|VSS \$1143 \$1322 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $818 r0 *1 28.055,1124.21 sg13_hv_nmos
M$818 \$1322 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $819 r0 *1 29.295,1124.21 sg13_hv_nmos
M$819 IOVSS|VSS \$1143 \$1323 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $820 r0 *1 31.075,1124.21 sg13_hv_nmos
M$820 \$1323 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $821 r0 *1 32.315,1124.21 sg13_hv_nmos
M$821 IOVSS|VSS \$1143 \$1324 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $822 r0 *1 34.095,1124.21 sg13_hv_nmos
M$822 \$1324 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $823 r0 *1 35.335,1124.21 sg13_hv_nmos
M$823 IOVSS|VSS \$1143 \$1325 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $824 r0 *1 37.115,1124.21 sg13_hv_nmos
M$824 \$1325 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $825 r0 *1 38.355,1124.21 sg13_hv_nmos
M$825 IOVSS|VSS \$1143 \$1326 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $826 r0 *1 40.135,1124.21 sg13_hv_nmos
M$826 \$1326 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $827 r0 *1 41.375,1124.21 sg13_hv_nmos
M$827 IOVSS|VSS \$1143 \$1327 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $828 r0 *1 43.155,1124.21 sg13_hv_nmos
M$828 \$1327 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $829 r0 *1 44.395,1124.21 sg13_hv_nmos
M$829 IOVSS|VSS \$1143 \$1328 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $830 r0 *1 46.175,1124.21 sg13_hv_nmos
M$830 \$1328 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $831 r0 *1 47.415,1124.21 sg13_hv_nmos
M$831 IOVSS|VSS \$1143 \$1329 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $832 r0 *1 49.195,1124.21 sg13_hv_nmos
M$832 \$1329 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $833 r0 *1 50.435,1124.21 sg13_hv_nmos
M$833 IOVSS|VSS \$1143 \$1330 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $834 r0 *1 52.215,1124.21 sg13_hv_nmos
M$834 \$1330 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $835 r0 *1 53.455,1124.21 sg13_hv_nmos
M$835 IOVSS|VSS \$1143 \$1331 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $836 r0 *1 55.235,1124.21 sg13_hv_nmos
M$836 \$1331 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $837 r0 *1 56.475,1124.21 sg13_hv_nmos
M$837 IOVSS|VSS \$1143 \$1332 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $838 r0 *1 58.255,1124.21 sg13_hv_nmos
M$838 \$1332 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $839 r0 *1 59.495,1124.21 sg13_hv_nmos
M$839 IOVSS|VSS \$1143 \$1333 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $840 r0 *1 61.275,1124.21 sg13_hv_nmos
M$840 \$1333 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $841 r0 *1 62.515,1124.21 sg13_hv_nmos
M$841 IOVSS|VSS \$1143 \$1334 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $842 r0 *1 64.295,1124.21 sg13_hv_nmos
M$842 \$1334 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $843 r0 *1 65.535,1124.21 sg13_hv_nmos
M$843 IOVSS|VSS \$1143 \$1335 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $844 r0 *1 67.315,1124.21 sg13_hv_nmos
M$844 \$1335 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $845 r0 *1 68.555,1124.21 sg13_hv_nmos
M$845 IOVSS|VSS \$1143 \$1336 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $846 r0 *1 70.335,1124.21 sg13_hv_nmos
M$846 \$1336 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $847 r0 *1 71.575,1124.21 sg13_hv_nmos
M$847 IOVSS|VSS \$1143 \$1337 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $848 r0 *1 308.155,1124.21 sg13_hv_nmos
M$848 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $849 r0 *1 309.935,1124.21 sg13_hv_nmos
M$849 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $850 r0 *1 311.175,1124.21 sg13_hv_nmos
M$850 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $851 r0 *1 312.955,1124.21 sg13_hv_nmos
M$851 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $852 r0 *1 314.195,1124.21 sg13_hv_nmos
M$852 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $853 r0 *1 315.975,1124.21 sg13_hv_nmos
M$853 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $854 r0 *1 317.215,1124.21 sg13_hv_nmos
M$854 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $855 r0 *1 318.995,1124.21 sg13_hv_nmos
M$855 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $856 r0 *1 320.235,1124.21 sg13_hv_nmos
M$856 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $857 r0 *1 322.015,1124.21 sg13_hv_nmos
M$857 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $858 r0 *1 323.255,1124.21 sg13_hv_nmos
M$858 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $859 r0 *1 325.035,1124.21 sg13_hv_nmos
M$859 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $860 r0 *1 326.275,1124.21 sg13_hv_nmos
M$860 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $861 r0 *1 328.055,1124.21 sg13_hv_nmos
M$861 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $862 r0 *1 329.295,1124.21 sg13_hv_nmos
M$862 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $863 r0 *1 331.075,1124.21 sg13_hv_nmos
M$863 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $864 r0 *1 332.315,1124.21 sg13_hv_nmos
M$864 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $865 r0 *1 334.095,1124.21 sg13_hv_nmos
M$865 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $866 r0 *1 335.335,1124.21 sg13_hv_nmos
M$866 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $867 r0 *1 337.115,1124.21 sg13_hv_nmos
M$867 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $868 r0 *1 338.355,1124.21 sg13_hv_nmos
M$868 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $869 r0 *1 340.135,1124.21 sg13_hv_nmos
M$869 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $870 r0 *1 341.375,1124.21 sg13_hv_nmos
M$870 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $871 r0 *1 343.155,1124.21 sg13_hv_nmos
M$871 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $872 r0 *1 344.395,1124.21 sg13_hv_nmos
M$872 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $873 r0 *1 346.175,1124.21 sg13_hv_nmos
M$873 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $874 r0 *1 347.415,1124.21 sg13_hv_nmos
M$874 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $875 r0 *1 349.195,1124.21 sg13_hv_nmos
M$875 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $876 r0 *1 350.435,1124.21 sg13_hv_nmos
M$876 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $877 r0 *1 352.215,1124.21 sg13_hv_nmos
M$877 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $878 r0 *1 353.455,1124.21 sg13_hv_nmos
M$878 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $879 r0 *1 355.235,1124.21 sg13_hv_nmos
M$879 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $880 r0 *1 356.475,1124.21 sg13_hv_nmos
M$880 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $881 r0 *1 358.255,1124.21 sg13_hv_nmos
M$881 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $882 r0 *1 359.495,1124.21 sg13_hv_nmos
M$882 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $883 r0 *1 361.275,1124.21 sg13_hv_nmos
M$883 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $884 r0 *1 362.515,1124.21 sg13_hv_nmos
M$884 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $885 r0 *1 364.295,1124.21 sg13_hv_nmos
M$885 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $886 r0 *1 365.535,1124.21 sg13_hv_nmos
M$886 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $887 r0 *1 367.315,1124.21 sg13_hv_nmos
M$887 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $888 r0 *1 368.555,1124.21 sg13_hv_nmos
M$888 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $889 r0 *1 370.335,1124.21 sg13_hv_nmos
M$889 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $890 r0 *1 371.575,1124.21 sg13_hv_nmos
M$890 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $891 r0 *1 708.155,1124.21 sg13_hv_nmos
M$891 IOVSS|VSS \$1145 \$1338 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $892 r0 *1 709.935,1124.21 sg13_hv_nmos
M$892 \$1338 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $893 r0 *1 711.175,1124.21 sg13_hv_nmos
M$893 IOVSS|VSS \$1145 \$1339 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $894 r0 *1 712.955,1124.21 sg13_hv_nmos
M$894 \$1339 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $895 r0 *1 714.195,1124.21 sg13_hv_nmos
M$895 IOVSS|VSS \$1145 \$1340 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $896 r0 *1 715.975,1124.21 sg13_hv_nmos
M$896 \$1340 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $897 r0 *1 717.215,1124.21 sg13_hv_nmos
M$897 IOVSS|VSS \$1145 \$1341 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $898 r0 *1 718.995,1124.21 sg13_hv_nmos
M$898 \$1341 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $899 r0 *1 720.235,1124.21 sg13_hv_nmos
M$899 IOVSS|VSS \$1145 \$1342 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $900 r0 *1 722.015,1124.21 sg13_hv_nmos
M$900 \$1342 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $901 r0 *1 723.255,1124.21 sg13_hv_nmos
M$901 IOVSS|VSS \$1145 \$1343 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $902 r0 *1 725.035,1124.21 sg13_hv_nmos
M$902 \$1343 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $903 r0 *1 726.275,1124.21 sg13_hv_nmos
M$903 IOVSS|VSS \$1145 \$1344 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $904 r0 *1 728.055,1124.21 sg13_hv_nmos
M$904 \$1344 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $905 r0 *1 729.295,1124.21 sg13_hv_nmos
M$905 IOVSS|VSS \$1145 \$1345 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $906 r0 *1 731.075,1124.21 sg13_hv_nmos
M$906 \$1345 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $907 r0 *1 732.315,1124.21 sg13_hv_nmos
M$907 IOVSS|VSS \$1145 \$1346 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $908 r0 *1 734.095,1124.21 sg13_hv_nmos
M$908 \$1346 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $909 r0 *1 735.335,1124.21 sg13_hv_nmos
M$909 IOVSS|VSS \$1145 \$1347 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $910 r0 *1 737.115,1124.21 sg13_hv_nmos
M$910 \$1347 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $911 r0 *1 738.355,1124.21 sg13_hv_nmos
M$911 IOVSS|VSS \$1145 \$1348 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $912 r0 *1 740.135,1124.21 sg13_hv_nmos
M$912 \$1348 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $913 r0 *1 741.375,1124.21 sg13_hv_nmos
M$913 IOVSS|VSS \$1145 \$1349 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $914 r0 *1 743.155,1124.21 sg13_hv_nmos
M$914 \$1349 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $915 r0 *1 744.395,1124.21 sg13_hv_nmos
M$915 IOVSS|VSS \$1145 \$1350 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $916 r0 *1 746.175,1124.21 sg13_hv_nmos
M$916 \$1350 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $917 r0 *1 747.415,1124.21 sg13_hv_nmos
M$917 IOVSS|VSS \$1145 \$1351 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $918 r0 *1 749.195,1124.21 sg13_hv_nmos
M$918 \$1351 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $919 r0 *1 750.435,1124.21 sg13_hv_nmos
M$919 IOVSS|VSS \$1145 \$1352 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $920 r0 *1 752.215,1124.21 sg13_hv_nmos
M$920 \$1352 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $921 r0 *1 753.455,1124.21 sg13_hv_nmos
M$921 IOVSS|VSS \$1145 \$1353 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $922 r0 *1 755.235,1124.21 sg13_hv_nmos
M$922 \$1353 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $923 r0 *1 756.475,1124.21 sg13_hv_nmos
M$923 IOVSS|VSS \$1145 \$1354 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $924 r0 *1 758.255,1124.21 sg13_hv_nmos
M$924 \$1354 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $925 r0 *1 759.495,1124.21 sg13_hv_nmos
M$925 IOVSS|VSS \$1145 \$1355 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $926 r0 *1 761.275,1124.21 sg13_hv_nmos
M$926 \$1355 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $927 r0 *1 762.515,1124.21 sg13_hv_nmos
M$927 IOVSS|VSS \$1145 \$1356 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $928 r0 *1 764.295,1124.21 sg13_hv_nmos
M$928 \$1356 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $929 r0 *1 765.535,1124.21 sg13_hv_nmos
M$929 IOVSS|VSS \$1145 \$1357 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $930 r0 *1 767.315,1124.21 sg13_hv_nmos
M$930 \$1357 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $931 r0 *1 768.555,1124.21 sg13_hv_nmos
M$931 IOVSS|VSS \$1145 \$1358 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $932 r0 *1 770.335,1124.21 sg13_hv_nmos
M$932 \$1358 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $933 r0 *1 771.575,1124.21 sg13_hv_nmos
M$933 IOVSS|VSS \$1145 \$1359 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $934 r0 *1 8.155,1129.05 sg13_hv_nmos
M$934 IOVSS|VSS \$1143 \$1316 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $935 r0 *1 9.935,1129.05 sg13_hv_nmos
M$935 \$1316 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $936 r0 *1 11.175,1129.05 sg13_hv_nmos
M$936 IOVSS|VSS \$1143 \$1317 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $937 r0 *1 12.955,1129.05 sg13_hv_nmos
M$937 \$1317 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $938 r0 *1 14.195,1129.05 sg13_hv_nmos
M$938 IOVSS|VSS \$1143 \$1318 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $939 r0 *1 15.975,1129.05 sg13_hv_nmos
M$939 \$1318 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $940 r0 *1 17.215,1129.05 sg13_hv_nmos
M$940 IOVSS|VSS \$1143 \$1319 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $941 r0 *1 18.995,1129.05 sg13_hv_nmos
M$941 \$1319 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $942 r0 *1 20.235,1129.05 sg13_hv_nmos
M$942 IOVSS|VSS \$1143 \$1320 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $943 r0 *1 22.015,1129.05 sg13_hv_nmos
M$943 \$1320 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $944 r0 *1 23.255,1129.05 sg13_hv_nmos
M$944 IOVSS|VSS \$1143 \$1321 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $945 r0 *1 25.035,1129.05 sg13_hv_nmos
M$945 \$1321 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $946 r0 *1 26.275,1129.05 sg13_hv_nmos
M$946 IOVSS|VSS \$1143 \$1322 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $947 r0 *1 28.055,1129.05 sg13_hv_nmos
M$947 \$1322 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $948 r0 *1 29.295,1129.05 sg13_hv_nmos
M$948 IOVSS|VSS \$1143 \$1323 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $949 r0 *1 31.075,1129.05 sg13_hv_nmos
M$949 \$1323 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $950 r0 *1 32.315,1129.05 sg13_hv_nmos
M$950 IOVSS|VSS \$1143 \$1324 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $951 r0 *1 34.095,1129.05 sg13_hv_nmos
M$951 \$1324 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $952 r0 *1 35.335,1129.05 sg13_hv_nmos
M$952 IOVSS|VSS \$1143 \$1325 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $953 r0 *1 37.115,1129.05 sg13_hv_nmos
M$953 \$1325 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $954 r0 *1 38.355,1129.05 sg13_hv_nmos
M$954 IOVSS|VSS \$1143 \$1326 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $955 r0 *1 40.135,1129.05 sg13_hv_nmos
M$955 \$1326 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $956 r0 *1 41.375,1129.05 sg13_hv_nmos
M$956 IOVSS|VSS \$1143 \$1327 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $957 r0 *1 43.155,1129.05 sg13_hv_nmos
M$957 \$1327 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $958 r0 *1 44.395,1129.05 sg13_hv_nmos
M$958 IOVSS|VSS \$1143 \$1328 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $959 r0 *1 46.175,1129.05 sg13_hv_nmos
M$959 \$1328 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $960 r0 *1 47.415,1129.05 sg13_hv_nmos
M$960 IOVSS|VSS \$1143 \$1329 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $961 r0 *1 49.195,1129.05 sg13_hv_nmos
M$961 \$1329 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $962 r0 *1 50.435,1129.05 sg13_hv_nmos
M$962 IOVSS|VSS \$1143 \$1330 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $963 r0 *1 52.215,1129.05 sg13_hv_nmos
M$963 \$1330 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $964 r0 *1 53.455,1129.05 sg13_hv_nmos
M$964 IOVSS|VSS \$1143 \$1331 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $965 r0 *1 55.235,1129.05 sg13_hv_nmos
M$965 \$1331 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $966 r0 *1 56.475,1129.05 sg13_hv_nmos
M$966 IOVSS|VSS \$1143 \$1332 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $967 r0 *1 58.255,1129.05 sg13_hv_nmos
M$967 \$1332 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $968 r0 *1 59.495,1129.05 sg13_hv_nmos
M$968 IOVSS|VSS \$1143 \$1333 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $969 r0 *1 61.275,1129.05 sg13_hv_nmos
M$969 \$1333 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $970 r0 *1 62.515,1129.05 sg13_hv_nmos
M$970 IOVSS|VSS \$1143 \$1334 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $971 r0 *1 64.295,1129.05 sg13_hv_nmos
M$971 \$1334 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $972 r0 *1 65.535,1129.05 sg13_hv_nmos
M$972 IOVSS|VSS \$1143 \$1335 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $973 r0 *1 67.315,1129.05 sg13_hv_nmos
M$973 \$1335 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $974 r0 *1 68.555,1129.05 sg13_hv_nmos
M$974 IOVSS|VSS \$1143 \$1336 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $975 r0 *1 70.335,1129.05 sg13_hv_nmos
M$975 \$1336 \$1143 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $976 r0 *1 71.575,1129.05 sg13_hv_nmos
M$976 IOVSS|VSS \$1143 \$1337 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $977 r0 *1 125.52,1129.05 sg13_hv_nmos
M$977 IOVSS|VSS \$1397 PAD|VREF IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $978 r0 *1 127.3,1129.05 sg13_hv_nmos
M$978 PAD|VREF \$1397 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $979 r0 *1 128.54,1129.05 sg13_hv_nmos
M$979 IOVSS|VSS \$1397 PAD|VREF IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $980 r0 *1 130.32,1129.05 sg13_hv_nmos
M$980 PAD|VREF \$1397 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $981 r0 *1 131.56,1129.05 sg13_hv_nmos
M$981 IOVSS|VSS \$1397 PAD|VREF IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $982 r0 *1 133.34,1129.05 sg13_hv_nmos
M$982 PAD|VREF \$1397 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $983 r0 *1 134.58,1129.05 sg13_hv_nmos
M$983 IOVSS|VSS \$1397 PAD|VREF IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $984 r0 *1 136.36,1129.05 sg13_hv_nmos
M$984 PAD|VREF \$1397 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $985 r0 *1 137.6,1129.05 sg13_hv_nmos
M$985 IOVSS|VSS \$1397 PAD|VREF IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $986 r0 *1 139.38,1129.05 sg13_hv_nmos
M$986 PAD|VREF \$1397 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $987 r0 *1 140.62,1129.05 sg13_hv_nmos
M$987 IOVSS|VSS \$1397 PAD|VREF IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $988 r0 *1 142.4,1129.05 sg13_hv_nmos
M$988 PAD|VREF \$1397 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $989 r0 *1 143.64,1129.05 sg13_hv_nmos
M$989 IOVSS|VSS \$1397 PAD|VREF IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $990 r0 *1 145.42,1129.05 sg13_hv_nmos
M$990 PAD|VREF \$1397 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $991 r0 *1 146.66,1129.05 sg13_hv_nmos
M$991 IOVSS|VSS \$1397 PAD|VREF IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $992 r0 *1 148.44,1129.05 sg13_hv_nmos
M$992 PAD|VREF \$1397 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $993 r0 *1 149.68,1129.05 sg13_hv_nmos
M$993 IOVSS|VSS \$1397 PAD|VREF IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $994 r0 *1 151.46,1129.05 sg13_hv_nmos
M$994 PAD|VREF \$1397 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $995 r0 *1 152.7,1129.05 sg13_hv_nmos
M$995 IOVSS|VSS \$1397 PAD|VREF IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $996 r0 *1 154.48,1129.05 sg13_hv_nmos
M$996 PAD|VREF \$1397 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $997 r0 *1 225.52,1129.05 sg13_hv_nmos
M$997 IOVSS|VSS \$1398 PAD|VLDO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $998 r0 *1 227.3,1129.05 sg13_hv_nmos
M$998 PAD|VLDO \$1398 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $999 r0 *1 228.54,1129.05 sg13_hv_nmos
M$999 IOVSS|VSS \$1398 PAD|VLDO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1000 r0 *1 230.32,1129.05 sg13_hv_nmos
M$1000 PAD|VLDO \$1398 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1001 r0 *1 231.56,1129.05 sg13_hv_nmos
M$1001 IOVSS|VSS \$1398 PAD|VLDO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1002 r0 *1 233.34,1129.05 sg13_hv_nmos
M$1002 PAD|VLDO \$1398 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1003 r0 *1 234.58,1129.05 sg13_hv_nmos
M$1003 IOVSS|VSS \$1398 PAD|VLDO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1004 r0 *1 236.36,1129.05 sg13_hv_nmos
M$1004 PAD|VLDO \$1398 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1005 r0 *1 237.6,1129.05 sg13_hv_nmos
M$1005 IOVSS|VSS \$1398 PAD|VLDO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1006 r0 *1 239.38,1129.05 sg13_hv_nmos
M$1006 PAD|VLDO \$1398 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1007 r0 *1 240.62,1129.05 sg13_hv_nmos
M$1007 IOVSS|VSS \$1398 PAD|VLDO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1008 r0 *1 242.4,1129.05 sg13_hv_nmos
M$1008 PAD|VLDO \$1398 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1009 r0 *1 243.64,1129.05 sg13_hv_nmos
M$1009 IOVSS|VSS \$1398 PAD|VLDO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1010 r0 *1 245.42,1129.05 sg13_hv_nmos
M$1010 PAD|VLDO \$1398 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1011 r0 *1 246.66,1129.05 sg13_hv_nmos
M$1011 IOVSS|VSS \$1398 PAD|VLDO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1012 r0 *1 248.44,1129.05 sg13_hv_nmos
M$1012 PAD|VLDO \$1398 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1013 r0 *1 249.68,1129.05 sg13_hv_nmos
M$1013 IOVSS|VSS \$1398 PAD|VLDO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1014 r0 *1 251.46,1129.05 sg13_hv_nmos
M$1014 PAD|VLDO \$1398 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1015 r0 *1 252.7,1129.05 sg13_hv_nmos
M$1015 IOVSS|VSS \$1398 PAD|VLDO IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1016 r0 *1 254.48,1129.05 sg13_hv_nmos
M$1016 PAD|VLDO \$1398 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1017 r0 *1 308.155,1129.05 sg13_hv_nmos
M$1017 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1018 r0 *1 309.935,1129.05 sg13_hv_nmos
M$1018 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1019 r0 *1 311.175,1129.05 sg13_hv_nmos
M$1019 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1020 r0 *1 312.955,1129.05 sg13_hv_nmos
M$1020 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1021 r0 *1 314.195,1129.05 sg13_hv_nmos
M$1021 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1022 r0 *1 315.975,1129.05 sg13_hv_nmos
M$1022 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1023 r0 *1 317.215,1129.05 sg13_hv_nmos
M$1023 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1024 r0 *1 318.995,1129.05 sg13_hv_nmos
M$1024 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1025 r0 *1 320.235,1129.05 sg13_hv_nmos
M$1025 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1026 r0 *1 322.015,1129.05 sg13_hv_nmos
M$1026 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1027 r0 *1 323.255,1129.05 sg13_hv_nmos
M$1027 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1028 r0 *1 325.035,1129.05 sg13_hv_nmos
M$1028 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1029 r0 *1 326.275,1129.05 sg13_hv_nmos
M$1029 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1030 r0 *1 328.055,1129.05 sg13_hv_nmos
M$1030 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1031 r0 *1 329.295,1129.05 sg13_hv_nmos
M$1031 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1032 r0 *1 331.075,1129.05 sg13_hv_nmos
M$1032 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1033 r0 *1 332.315,1129.05 sg13_hv_nmos
M$1033 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1034 r0 *1 334.095,1129.05 sg13_hv_nmos
M$1034 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1035 r0 *1 335.335,1129.05 sg13_hv_nmos
M$1035 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1036 r0 *1 337.115,1129.05 sg13_hv_nmos
M$1036 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1037 r0 *1 338.355,1129.05 sg13_hv_nmos
M$1037 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1038 r0 *1 340.135,1129.05 sg13_hv_nmos
M$1038 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1039 r0 *1 341.375,1129.05 sg13_hv_nmos
M$1039 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1040 r0 *1 343.155,1129.05 sg13_hv_nmos
M$1040 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1041 r0 *1 344.395,1129.05 sg13_hv_nmos
M$1041 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1042 r0 *1 346.175,1129.05 sg13_hv_nmos
M$1042 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1043 r0 *1 347.415,1129.05 sg13_hv_nmos
M$1043 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1044 r0 *1 349.195,1129.05 sg13_hv_nmos
M$1044 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1045 r0 *1 350.435,1129.05 sg13_hv_nmos
M$1045 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1046 r0 *1 352.215,1129.05 sg13_hv_nmos
M$1046 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1047 r0 *1 353.455,1129.05 sg13_hv_nmos
M$1047 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1048 r0 *1 355.235,1129.05 sg13_hv_nmos
M$1048 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1049 r0 *1 356.475,1129.05 sg13_hv_nmos
M$1049 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1050 r0 *1 358.255,1129.05 sg13_hv_nmos
M$1050 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1051 r0 *1 359.495,1129.05 sg13_hv_nmos
M$1051 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1052 r0 *1 361.275,1129.05 sg13_hv_nmos
M$1052 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1053 r0 *1 362.515,1129.05 sg13_hv_nmos
M$1053 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1054 r0 *1 364.295,1129.05 sg13_hv_nmos
M$1054 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1055 r0 *1 365.535,1129.05 sg13_hv_nmos
M$1055 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1056 r0 *1 367.315,1129.05 sg13_hv_nmos
M$1056 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1057 r0 *1 368.555,1129.05 sg13_hv_nmos
M$1057 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1058 r0 *1 370.335,1129.05 sg13_hv_nmos
M$1058 IOVDD \$1144 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1059 r0 *1 371.575,1129.05 sg13_hv_nmos
M$1059 IOVSS|VSS \$1144 IOVDD IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1060 r0 *1 708.155,1129.05 sg13_hv_nmos
M$1060 IOVSS|VSS \$1145 \$1338 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1061 r0 *1 709.935,1129.05 sg13_hv_nmos
M$1061 \$1338 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1062 r0 *1 711.175,1129.05 sg13_hv_nmos
M$1062 IOVSS|VSS \$1145 \$1339 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1063 r0 *1 712.955,1129.05 sg13_hv_nmos
M$1063 \$1339 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1064 r0 *1 714.195,1129.05 sg13_hv_nmos
M$1064 IOVSS|VSS \$1145 \$1340 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1065 r0 *1 715.975,1129.05 sg13_hv_nmos
M$1065 \$1340 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1066 r0 *1 717.215,1129.05 sg13_hv_nmos
M$1066 IOVSS|VSS \$1145 \$1341 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1067 r0 *1 718.995,1129.05 sg13_hv_nmos
M$1067 \$1341 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1068 r0 *1 720.235,1129.05 sg13_hv_nmos
M$1068 IOVSS|VSS \$1145 \$1342 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1069 r0 *1 722.015,1129.05 sg13_hv_nmos
M$1069 \$1342 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1070 r0 *1 723.255,1129.05 sg13_hv_nmos
M$1070 IOVSS|VSS \$1145 \$1343 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1071 r0 *1 725.035,1129.05 sg13_hv_nmos
M$1071 \$1343 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1072 r0 *1 726.275,1129.05 sg13_hv_nmos
M$1072 IOVSS|VSS \$1145 \$1344 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1073 r0 *1 728.055,1129.05 sg13_hv_nmos
M$1073 \$1344 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1074 r0 *1 729.295,1129.05 sg13_hv_nmos
M$1074 IOVSS|VSS \$1145 \$1345 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1075 r0 *1 731.075,1129.05 sg13_hv_nmos
M$1075 \$1345 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1076 r0 *1 732.315,1129.05 sg13_hv_nmos
M$1076 IOVSS|VSS \$1145 \$1346 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1077 r0 *1 734.095,1129.05 sg13_hv_nmos
M$1077 \$1346 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1078 r0 *1 735.335,1129.05 sg13_hv_nmos
M$1078 IOVSS|VSS \$1145 \$1347 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1079 r0 *1 737.115,1129.05 sg13_hv_nmos
M$1079 \$1347 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1080 r0 *1 738.355,1129.05 sg13_hv_nmos
M$1080 IOVSS|VSS \$1145 \$1348 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1081 r0 *1 740.135,1129.05 sg13_hv_nmos
M$1081 \$1348 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1082 r0 *1 741.375,1129.05 sg13_hv_nmos
M$1082 IOVSS|VSS \$1145 \$1349 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1083 r0 *1 743.155,1129.05 sg13_hv_nmos
M$1083 \$1349 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1084 r0 *1 744.395,1129.05 sg13_hv_nmos
M$1084 IOVSS|VSS \$1145 \$1350 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1085 r0 *1 746.175,1129.05 sg13_hv_nmos
M$1085 \$1350 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1086 r0 *1 747.415,1129.05 sg13_hv_nmos
M$1086 IOVSS|VSS \$1145 \$1351 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1087 r0 *1 749.195,1129.05 sg13_hv_nmos
M$1087 \$1351 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1088 r0 *1 750.435,1129.05 sg13_hv_nmos
M$1088 IOVSS|VSS \$1145 \$1352 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1089 r0 *1 752.215,1129.05 sg13_hv_nmos
M$1089 \$1352 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1090 r0 *1 753.455,1129.05 sg13_hv_nmos
M$1090 IOVSS|VSS \$1145 \$1353 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1091 r0 *1 755.235,1129.05 sg13_hv_nmos
M$1091 \$1353 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1092 r0 *1 756.475,1129.05 sg13_hv_nmos
M$1092 IOVSS|VSS \$1145 \$1354 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1093 r0 *1 758.255,1129.05 sg13_hv_nmos
M$1093 \$1354 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1094 r0 *1 759.495,1129.05 sg13_hv_nmos
M$1094 IOVSS|VSS \$1145 \$1355 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1095 r0 *1 761.275,1129.05 sg13_hv_nmos
M$1095 \$1355 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1096 r0 *1 762.515,1129.05 sg13_hv_nmos
M$1096 IOVSS|VSS \$1145 \$1356 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1097 r0 *1 764.295,1129.05 sg13_hv_nmos
M$1097 \$1356 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1098 r0 *1 765.535,1129.05 sg13_hv_nmos
M$1098 IOVSS|VSS \$1145 \$1357 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1099 r0 *1 767.315,1129.05 sg13_hv_nmos
M$1099 \$1357 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1100 r0 *1 768.555,1129.05 sg13_hv_nmos
M$1100 IOVSS|VSS \$1145 \$1358 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1101 r0 *1 770.335,1129.05 sg13_hv_nmos
M$1101 \$1358 \$1145 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1102 r0 *1 771.575,1129.05 sg13_hv_nmos
M$1102 IOVSS|VSS \$1145 \$1359 IOVSS|VSS sg13_hv_nmos W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1103 r0 *1 240.255,163.995 sg13_lv_pmos
M$1103 res_c \$186 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1104 r0 *1 440.255,163.995 sg13_lv_pmos
M$1104 ck4_c \$187 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1105 r0 *1 540.255,163.995 sg13_lv_pmos
M$1105 ck5_c \$188 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1106 r0 *1 640.255,163.995 sg13_lv_pmos
M$1106 ck6_c \$189 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1107 r0 *1 796.005,217.48 sg13_lv_pmos
M$1107 \$237 out6_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1108 r0 *1 796.005,220.99 sg13_lv_pmos
M$1108 \$264 out6_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1109 r0 *1 796.005,317.48 sg13_lv_pmos
M$1109 \$350 out5_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1110 r0 *1 796.005,320.99 sg13_lv_pmos
M$1110 \$377 out5_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1111 r0 *1 796.005,417.48 sg13_lv_pmos
M$1111 \$463 out4_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1112 r0 *1 796.005,420.99 sg13_lv_pmos
M$1112 \$490 out4_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1113 r0 *1 796.005,717.48 sg13_lv_pmos
M$1113 \$750 out3_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1114 r0 *1 796.005,720.99 sg13_lv_pmos
M$1114 \$777 out3_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1115 r0 *1 796.005,817.48 sg13_lv_pmos
M$1115 \$863 out2_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1116 r0 *1 796.005,820.99 sg13_lv_pmos
M$1116 \$890 out2_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1117 r0 *1 796.005,917.48 sg13_lv_pmos
M$1117 \$976 out1_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1118 r0 *1 796.005,920.99 sg13_lv_pmos
M$1118 \$1003 out1_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1119 r0 *1 440.255,976.005 sg13_lv_pmos
M$1119 ck3_c \$1067 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1120 r0 *1 540.255,976.005 sg13_lv_pmos
M$1120 ck2_c \$1068 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1121 r0 *1 640.255,976.005 sg13_lv_pmos
M$1121 ck1_c \$1069 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1122 r0 *1 241.765,163.945 sg13_hv_pmos
M$1122 VDD \$129 \$186 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1123 r0 *1 441.765,163.945 sg13_hv_pmos
M$1123 VDD \$130 \$187 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1124 r0 *1 541.765,163.945 sg13_hv_pmos
M$1124 VDD \$132 \$188 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1125 r0 *1 641.765,163.945 sg13_hv_pmos
M$1125 VDD \$133 \$189 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1126 r0 *1 -108.92,205.52 sg13_hv_pmos
M$1126 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1127 r0 *1 -108.92,207.3 sg13_hv_pmos
M$1127 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1128 r0 *1 -108.92,208.54 sg13_hv_pmos
M$1128 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1129 r0 *1 -108.92,210.32 sg13_hv_pmos
M$1129 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1130 r0 *1 -108.92,211.56 sg13_hv_pmos
M$1130 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1131 r0 *1 -108.92,213.34 sg13_hv_pmos
M$1131 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1132 r0 *1 -108.92,214.58 sg13_hv_pmos
M$1132 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1133 r0 *1 -108.92,216.36 sg13_hv_pmos
M$1133 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1134 r0 *1 -108.92,217.6 sg13_hv_pmos
M$1134 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1135 r0 *1 -108.92,219.38 sg13_hv_pmos
M$1135 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1136 r0 *1 -108.92,220.62 sg13_hv_pmos
M$1136 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1137 r0 *1 -108.92,222.4 sg13_hv_pmos
M$1137 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1138 r0 *1 -108.92,223.64 sg13_hv_pmos
M$1138 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1139 r0 *1 -108.92,225.42 sg13_hv_pmos
M$1139 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1140 r0 *1 -108.92,226.66 sg13_hv_pmos
M$1140 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1141 r0 *1 -108.92,228.44 sg13_hv_pmos
M$1141 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1142 r0 *1 -108.92,229.68 sg13_hv_pmos
M$1142 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1143 r0 *1 -108.92,231.46 sg13_hv_pmos
M$1143 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1144 r0 *1 -108.92,232.7 sg13_hv_pmos
M$1144 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1145 r0 *1 -108.92,234.48 sg13_hv_pmos
M$1145 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1146 r0 *1 -101.82,205.52 sg13_hv_pmos
M$1146 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1147 r0 *1 -101.82,207.3 sg13_hv_pmos
M$1147 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1148 r0 *1 -101.82,208.54 sg13_hv_pmos
M$1148 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1149 r0 *1 -101.82,210.32 sg13_hv_pmos
M$1149 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1150 r0 *1 -101.82,211.56 sg13_hv_pmos
M$1150 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1151 r0 *1 -101.82,213.34 sg13_hv_pmos
M$1151 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1152 r0 *1 -101.82,214.58 sg13_hv_pmos
M$1152 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1153 r0 *1 -101.82,216.36 sg13_hv_pmos
M$1153 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1154 r0 *1 -101.82,217.6 sg13_hv_pmos
M$1154 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1155 r0 *1 -101.82,219.38 sg13_hv_pmos
M$1155 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1156 r0 *1 -101.82,220.62 sg13_hv_pmos
M$1156 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1157 r0 *1 -101.82,222.4 sg13_hv_pmos
M$1157 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1158 r0 *1 -101.82,223.64 sg13_hv_pmos
M$1158 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1159 r0 *1 -101.82,225.42 sg13_hv_pmos
M$1159 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1160 r0 *1 -101.82,226.66 sg13_hv_pmos
M$1160 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1161 r0 *1 -101.82,228.44 sg13_hv_pmos
M$1161 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1162 r0 *1 -101.82,229.68 sg13_hv_pmos
M$1162 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1163 r0 *1 -101.82,231.46 sg13_hv_pmos
M$1163 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1164 r0 *1 -101.82,232.7 sg13_hv_pmos
M$1164 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1165 r0 *1 -101.82,234.48 sg13_hv_pmos
M$1165 IN6|PAD \$228 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1166 r0 *1 881.82,214.58 sg13_hv_pmos
M$1166 IOVDD \$218 OUT6 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1167 r0 *1 881.82,216.36 sg13_hv_pmos
M$1167 OUT6 \$218 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1168 r0 *1 881.82,217.6 sg13_hv_pmos
M$1168 IOVDD \$218 OUT6 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1169 r0 *1 881.82,219.38 sg13_hv_pmos
M$1169 OUT6 \$218 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1170 r0 *1 881.82,220.62 sg13_hv_pmos
M$1170 IOVDD \$218 OUT6 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1171 r0 *1 881.82,222.4 sg13_hv_pmos
M$1171 OUT6 \$218 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1172 r0 *1 881.82,223.64 sg13_hv_pmos
M$1172 IOVDD \$218 OUT6 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1173 r0 *1 881.82,225.42 sg13_hv_pmos
M$1173 OUT6 \$218 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1174 r0 *1 888.92,214.58 sg13_hv_pmos
M$1174 IOVDD \$218 OUT6 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1175 r0 *1 888.92,216.36 sg13_hv_pmos
M$1175 OUT6 \$218 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1176 r0 *1 888.92,217.6 sg13_hv_pmos
M$1176 IOVDD \$218 OUT6 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1177 r0 *1 888.92,219.38 sg13_hv_pmos
M$1177 OUT6 \$218 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1178 r0 *1 888.92,220.62 sg13_hv_pmos
M$1178 IOVDD \$218 OUT6 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1179 r0 *1 888.92,222.4 sg13_hv_pmos
M$1179 OUT6 \$218 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1180 r0 *1 888.92,223.64 sg13_hv_pmos
M$1180 IOVDD \$218 OUT6 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1181 r0 *1 888.92,225.42 sg13_hv_pmos
M$1181 OUT6 \$218 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1182 r0 *1 808.82,217.64 sg13_hv_pmos
M$1182 \$238 \$248 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1183 r0 *1 808.82,218.47 sg13_hv_pmos
M$1183 IOVDD \$238 \$248 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1184 r0 *1 808.82,219.81 sg13_hv_pmos
M$1184 IOVDD \$248 \$253 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1185 r0 *1 808.82,221.15 sg13_hv_pmos
M$1185 \$265 \$272 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1186 r0 *1 808.82,221.98 sg13_hv_pmos
M$1186 IOVDD \$265 \$272 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1187 r0 *1 808.82,223.32 sg13_hv_pmos
M$1187 IOVDD \$272 \$218 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1188 r0 *1 -108.92,305.52 sg13_hv_pmos
M$1188 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1189 r0 *1 -108.92,307.3 sg13_hv_pmos
M$1189 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1190 r0 *1 -108.92,308.54 sg13_hv_pmos
M$1190 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1191 r0 *1 -108.92,310.32 sg13_hv_pmos
M$1191 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1192 r0 *1 -108.92,311.56 sg13_hv_pmos
M$1192 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1193 r0 *1 -108.92,313.34 sg13_hv_pmos
M$1193 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1194 r0 *1 -108.92,314.58 sg13_hv_pmos
M$1194 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1195 r0 *1 -108.92,316.36 sg13_hv_pmos
M$1195 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1196 r0 *1 -108.92,317.6 sg13_hv_pmos
M$1196 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1197 r0 *1 -108.92,319.38 sg13_hv_pmos
M$1197 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1198 r0 *1 -108.92,320.62 sg13_hv_pmos
M$1198 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1199 r0 *1 -108.92,322.4 sg13_hv_pmos
M$1199 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1200 r0 *1 -108.92,323.64 sg13_hv_pmos
M$1200 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1201 r0 *1 -108.92,325.42 sg13_hv_pmos
M$1201 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1202 r0 *1 -108.92,326.66 sg13_hv_pmos
M$1202 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1203 r0 *1 -108.92,328.44 sg13_hv_pmos
M$1203 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1204 r0 *1 -108.92,329.68 sg13_hv_pmos
M$1204 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1205 r0 *1 -108.92,331.46 sg13_hv_pmos
M$1205 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1206 r0 *1 -108.92,332.7 sg13_hv_pmos
M$1206 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1207 r0 *1 -108.92,334.48 sg13_hv_pmos
M$1207 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1208 r0 *1 -101.82,305.52 sg13_hv_pmos
M$1208 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1209 r0 *1 -101.82,307.3 sg13_hv_pmos
M$1209 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1210 r0 *1 -101.82,308.54 sg13_hv_pmos
M$1210 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1211 r0 *1 -101.82,310.32 sg13_hv_pmos
M$1211 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1212 r0 *1 -101.82,311.56 sg13_hv_pmos
M$1212 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1213 r0 *1 -101.82,313.34 sg13_hv_pmos
M$1213 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1214 r0 *1 -101.82,314.58 sg13_hv_pmos
M$1214 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1215 r0 *1 -101.82,316.36 sg13_hv_pmos
M$1215 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1216 r0 *1 -101.82,317.6 sg13_hv_pmos
M$1216 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1217 r0 *1 -101.82,319.38 sg13_hv_pmos
M$1217 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1218 r0 *1 -101.82,320.62 sg13_hv_pmos
M$1218 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1219 r0 *1 -101.82,322.4 sg13_hv_pmos
M$1219 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1220 r0 *1 -101.82,323.64 sg13_hv_pmos
M$1220 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1221 r0 *1 -101.82,325.42 sg13_hv_pmos
M$1221 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1222 r0 *1 -101.82,326.66 sg13_hv_pmos
M$1222 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1223 r0 *1 -101.82,328.44 sg13_hv_pmos
M$1223 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1224 r0 *1 -101.82,329.68 sg13_hv_pmos
M$1224 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1225 r0 *1 -101.82,331.46 sg13_hv_pmos
M$1225 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1226 r0 *1 -101.82,332.7 sg13_hv_pmos
M$1226 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1227 r0 *1 -101.82,334.48 sg13_hv_pmos
M$1227 IN5|PAD \$341 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1228 r0 *1 881.82,314.58 sg13_hv_pmos
M$1228 IOVDD \$331 OUT5 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1229 r0 *1 881.82,316.36 sg13_hv_pmos
M$1229 OUT5 \$331 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1230 r0 *1 881.82,317.6 sg13_hv_pmos
M$1230 IOVDD \$331 OUT5 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1231 r0 *1 881.82,319.38 sg13_hv_pmos
M$1231 OUT5 \$331 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1232 r0 *1 881.82,320.62 sg13_hv_pmos
M$1232 IOVDD \$331 OUT5 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1233 r0 *1 881.82,322.4 sg13_hv_pmos
M$1233 OUT5 \$331 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1234 r0 *1 881.82,323.64 sg13_hv_pmos
M$1234 IOVDD \$331 OUT5 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1235 r0 *1 881.82,325.42 sg13_hv_pmos
M$1235 OUT5 \$331 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1236 r0 *1 888.92,314.58 sg13_hv_pmos
M$1236 IOVDD \$331 OUT5 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1237 r0 *1 888.92,316.36 sg13_hv_pmos
M$1237 OUT5 \$331 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1238 r0 *1 888.92,317.6 sg13_hv_pmos
M$1238 IOVDD \$331 OUT5 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1239 r0 *1 888.92,319.38 sg13_hv_pmos
M$1239 OUT5 \$331 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1240 r0 *1 888.92,320.62 sg13_hv_pmos
M$1240 IOVDD \$331 OUT5 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1241 r0 *1 888.92,322.4 sg13_hv_pmos
M$1241 OUT5 \$331 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1242 r0 *1 888.92,323.64 sg13_hv_pmos
M$1242 IOVDD \$331 OUT5 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1243 r0 *1 888.92,325.42 sg13_hv_pmos
M$1243 OUT5 \$331 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1244 r0 *1 808.82,317.64 sg13_hv_pmos
M$1244 \$351 \$361 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1245 r0 *1 808.82,318.47 sg13_hv_pmos
M$1245 IOVDD \$351 \$361 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1246 r0 *1 808.82,319.81 sg13_hv_pmos
M$1246 IOVDD \$361 \$366 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1247 r0 *1 808.82,321.15 sg13_hv_pmos
M$1247 \$378 \$385 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1248 r0 *1 808.82,321.98 sg13_hv_pmos
M$1248 IOVDD \$378 \$385 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1249 r0 *1 808.82,323.32 sg13_hv_pmos
M$1249 IOVDD \$385 \$331 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1250 r0 *1 -108.92,405.52 sg13_hv_pmos
M$1250 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1251 r0 *1 -108.92,407.3 sg13_hv_pmos
M$1251 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1252 r0 *1 -108.92,408.54 sg13_hv_pmos
M$1252 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1253 r0 *1 -108.92,410.32 sg13_hv_pmos
M$1253 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1254 r0 *1 -108.92,411.56 sg13_hv_pmos
M$1254 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1255 r0 *1 -108.92,413.34 sg13_hv_pmos
M$1255 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1256 r0 *1 -108.92,414.58 sg13_hv_pmos
M$1256 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1257 r0 *1 -108.92,416.36 sg13_hv_pmos
M$1257 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1258 r0 *1 -108.92,417.6 sg13_hv_pmos
M$1258 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1259 r0 *1 -108.92,419.38 sg13_hv_pmos
M$1259 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1260 r0 *1 -108.92,420.62 sg13_hv_pmos
M$1260 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1261 r0 *1 -108.92,422.4 sg13_hv_pmos
M$1261 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1262 r0 *1 -108.92,423.64 sg13_hv_pmos
M$1262 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1263 r0 *1 -108.92,425.42 sg13_hv_pmos
M$1263 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1264 r0 *1 -108.92,426.66 sg13_hv_pmos
M$1264 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1265 r0 *1 -108.92,428.44 sg13_hv_pmos
M$1265 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1266 r0 *1 -108.92,429.68 sg13_hv_pmos
M$1266 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1267 r0 *1 -108.92,431.46 sg13_hv_pmos
M$1267 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1268 r0 *1 -108.92,432.7 sg13_hv_pmos
M$1268 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1269 r0 *1 -108.92,434.48 sg13_hv_pmos
M$1269 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1270 r0 *1 -101.82,405.52 sg13_hv_pmos
M$1270 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1271 r0 *1 -101.82,407.3 sg13_hv_pmos
M$1271 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1272 r0 *1 -101.82,408.54 sg13_hv_pmos
M$1272 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1273 r0 *1 -101.82,410.32 sg13_hv_pmos
M$1273 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1274 r0 *1 -101.82,411.56 sg13_hv_pmos
M$1274 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1275 r0 *1 -101.82,413.34 sg13_hv_pmos
M$1275 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1276 r0 *1 -101.82,414.58 sg13_hv_pmos
M$1276 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1277 r0 *1 -101.82,416.36 sg13_hv_pmos
M$1277 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1278 r0 *1 -101.82,417.6 sg13_hv_pmos
M$1278 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1279 r0 *1 -101.82,419.38 sg13_hv_pmos
M$1279 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1280 r0 *1 -101.82,420.62 sg13_hv_pmos
M$1280 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1281 r0 *1 -101.82,422.4 sg13_hv_pmos
M$1281 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1282 r0 *1 -101.82,423.64 sg13_hv_pmos
M$1282 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1283 r0 *1 -101.82,425.42 sg13_hv_pmos
M$1283 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1284 r0 *1 -101.82,426.66 sg13_hv_pmos
M$1284 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1285 r0 *1 -101.82,428.44 sg13_hv_pmos
M$1285 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1286 r0 *1 -101.82,429.68 sg13_hv_pmos
M$1286 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1287 r0 *1 -101.82,431.46 sg13_hv_pmos
M$1287 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1288 r0 *1 -101.82,432.7 sg13_hv_pmos
M$1288 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1289 r0 *1 -101.82,434.48 sg13_hv_pmos
M$1289 IN4|PAD \$454 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1290 r0 *1 881.82,414.58 sg13_hv_pmos
M$1290 IOVDD \$444 OUT4 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1291 r0 *1 881.82,416.36 sg13_hv_pmos
M$1291 OUT4 \$444 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1292 r0 *1 881.82,417.6 sg13_hv_pmos
M$1292 IOVDD \$444 OUT4 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1293 r0 *1 881.82,419.38 sg13_hv_pmos
M$1293 OUT4 \$444 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1294 r0 *1 881.82,420.62 sg13_hv_pmos
M$1294 IOVDD \$444 OUT4 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1295 r0 *1 881.82,422.4 sg13_hv_pmos
M$1295 OUT4 \$444 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1296 r0 *1 881.82,423.64 sg13_hv_pmos
M$1296 IOVDD \$444 OUT4 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1297 r0 *1 881.82,425.42 sg13_hv_pmos
M$1297 OUT4 \$444 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1298 r0 *1 888.92,414.58 sg13_hv_pmos
M$1298 IOVDD \$444 OUT4 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1299 r0 *1 888.92,416.36 sg13_hv_pmos
M$1299 OUT4 \$444 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1300 r0 *1 888.92,417.6 sg13_hv_pmos
M$1300 IOVDD \$444 OUT4 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1301 r0 *1 888.92,419.38 sg13_hv_pmos
M$1301 OUT4 \$444 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1302 r0 *1 888.92,420.62 sg13_hv_pmos
M$1302 IOVDD \$444 OUT4 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1303 r0 *1 888.92,422.4 sg13_hv_pmos
M$1303 OUT4 \$444 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1304 r0 *1 888.92,423.64 sg13_hv_pmos
M$1304 IOVDD \$444 OUT4 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1305 r0 *1 888.92,425.42 sg13_hv_pmos
M$1305 OUT4 \$444 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1306 r0 *1 808.82,417.64 sg13_hv_pmos
M$1306 \$464 \$474 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1307 r0 *1 808.82,418.47 sg13_hv_pmos
M$1307 IOVDD \$464 \$474 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1308 r0 *1 808.82,419.81 sg13_hv_pmos
M$1308 IOVDD \$474 \$479 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1309 r0 *1 808.82,421.15 sg13_hv_pmos
M$1309 \$491 \$498 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1310 r0 *1 808.82,421.98 sg13_hv_pmos
M$1310 IOVDD \$491 \$498 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1311 r0 *1 808.82,423.32 sg13_hv_pmos
M$1311 IOVDD \$498 \$444 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1312 r0 *1 -108.92,505.52 sg13_hv_pmos
M$1312 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1313 r0 *1 -108.92,507.3 sg13_hv_pmos
M$1313 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1314 r0 *1 -108.92,508.54 sg13_hv_pmos
M$1314 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1315 r0 *1 -108.92,510.32 sg13_hv_pmos
M$1315 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1316 r0 *1 -108.92,511.56 sg13_hv_pmos
M$1316 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1317 r0 *1 -108.92,513.34 sg13_hv_pmos
M$1317 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1318 r0 *1 -108.92,514.58 sg13_hv_pmos
M$1318 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1319 r0 *1 -108.92,516.36 sg13_hv_pmos
M$1319 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1320 r0 *1 -108.92,517.6 sg13_hv_pmos
M$1320 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1321 r0 *1 -108.92,519.38 sg13_hv_pmos
M$1321 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1322 r0 *1 -108.92,520.62 sg13_hv_pmos
M$1322 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1323 r0 *1 -108.92,522.4 sg13_hv_pmos
M$1323 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1324 r0 *1 -108.92,523.64 sg13_hv_pmos
M$1324 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1325 r0 *1 -108.92,525.42 sg13_hv_pmos
M$1325 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1326 r0 *1 -108.92,526.66 sg13_hv_pmos
M$1326 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1327 r0 *1 -108.92,528.44 sg13_hv_pmos
M$1327 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1328 r0 *1 -108.92,529.68 sg13_hv_pmos
M$1328 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1329 r0 *1 -108.92,531.46 sg13_hv_pmos
M$1329 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1330 r0 *1 -108.92,532.7 sg13_hv_pmos
M$1330 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1331 r0 *1 -108.92,534.48 sg13_hv_pmos
M$1331 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1332 r0 *1 -101.82,505.52 sg13_hv_pmos
M$1332 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1333 r0 *1 -101.82,507.3 sg13_hv_pmos
M$1333 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1334 r0 *1 -101.82,508.54 sg13_hv_pmos
M$1334 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1335 r0 *1 -101.82,510.32 sg13_hv_pmos
M$1335 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1336 r0 *1 -101.82,511.56 sg13_hv_pmos
M$1336 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1337 r0 *1 -101.82,513.34 sg13_hv_pmos
M$1337 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1338 r0 *1 -101.82,514.58 sg13_hv_pmos
M$1338 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1339 r0 *1 -101.82,516.36 sg13_hv_pmos
M$1339 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1340 r0 *1 -101.82,517.6 sg13_hv_pmos
M$1340 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1341 r0 *1 -101.82,519.38 sg13_hv_pmos
M$1341 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1342 r0 *1 -101.82,520.62 sg13_hv_pmos
M$1342 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1343 r0 *1 -101.82,522.4 sg13_hv_pmos
M$1343 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1344 r0 *1 -101.82,523.64 sg13_hv_pmos
M$1344 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1345 r0 *1 -101.82,525.42 sg13_hv_pmos
M$1345 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1346 r0 *1 -101.82,526.66 sg13_hv_pmos
M$1346 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1347 r0 *1 -101.82,528.44 sg13_hv_pmos
M$1347 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1348 r0 *1 -101.82,529.68 sg13_hv_pmos
M$1348 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1349 r0 *1 -101.82,531.46 sg13_hv_pmos
M$1349 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1350 r0 *1 -101.82,532.7 sg13_hv_pmos
M$1350 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1351 r0 *1 -101.82,534.48 sg13_hv_pmos
M$1351 PAD|VLO \$569 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1352 r0 *1 865.09,598.44 sg13_hv_pmos
M$1352 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1353 r0 *1 865.09,599.32 sg13_hv_pmos
M$1353 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1354 r0 *1 865.09,600.2 sg13_hv_pmos
M$1354 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1355 r0 *1 865.09,601.08 sg13_hv_pmos
M$1355 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1356 r0 *1 865.09,601.96 sg13_hv_pmos
M$1356 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1357 r0 *1 865.09,602.84 sg13_hv_pmos
M$1357 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1358 r0 *1 865.09,603.72 sg13_hv_pmos
M$1358 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1359 r0 *1 865.09,604.6 sg13_hv_pmos
M$1359 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1360 r0 *1 865.09,605.48 sg13_hv_pmos
M$1360 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1361 r0 *1 865.09,606.36 sg13_hv_pmos
M$1361 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1362 r0 *1 865.09,607.24 sg13_hv_pmos
M$1362 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1363 r0 *1 865.09,608.12 sg13_hv_pmos
M$1363 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1364 r0 *1 865.09,609 sg13_hv_pmos
M$1364 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1365 r0 *1 865.09,609.88 sg13_hv_pmos
M$1365 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1366 r0 *1 865.09,610.76 sg13_hv_pmos
M$1366 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1367 r0 *1 865.09,611.64 sg13_hv_pmos
M$1367 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1368 r0 *1 865.09,612.52 sg13_hv_pmos
M$1368 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1369 r0 *1 865.09,613.4 sg13_hv_pmos
M$1369 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1370 r0 *1 865.09,614.28 sg13_hv_pmos
M$1370 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1371 r0 *1 865.09,615.16 sg13_hv_pmos
M$1371 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1372 r0 *1 865.09,616.04 sg13_hv_pmos
M$1372 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1373 r0 *1 865.09,616.92 sg13_hv_pmos
M$1373 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1374 r0 *1 865.09,617.8 sg13_hv_pmos
M$1374 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1375 r0 *1 865.09,618.68 sg13_hv_pmos
M$1375 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1376 r0 *1 865.09,619.56 sg13_hv_pmos
M$1376 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1377 r0 *1 865.09,620.44 sg13_hv_pmos
M$1377 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1378 r0 *1 865.09,621.32 sg13_hv_pmos
M$1378 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1379 r0 *1 865.09,622.2 sg13_hv_pmos
M$1379 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1380 r0 *1 865.09,623.08 sg13_hv_pmos
M$1380 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1381 r0 *1 865.09,623.96 sg13_hv_pmos
M$1381 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1382 r0 *1 865.09,624.84 sg13_hv_pmos
M$1382 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1383 r0 *1 865.09,625.72 sg13_hv_pmos
M$1383 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1384 r0 *1 865.09,626.6 sg13_hv_pmos
M$1384 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1385 r0 *1 865.09,627.48 sg13_hv_pmos
M$1385 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1386 r0 *1 865.09,628.36 sg13_hv_pmos
M$1386 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1387 r0 *1 865.09,629.24 sg13_hv_pmos
M$1387 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1388 r0 *1 865.09,630.12 sg13_hv_pmos
M$1388 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1389 r0 *1 865.09,631 sg13_hv_pmos
M$1389 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1390 r0 *1 865.09,631.88 sg13_hv_pmos
M$1390 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1391 r0 *1 865.09,632.76 sg13_hv_pmos
M$1391 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1392 r0 *1 865.09,633.64 sg13_hv_pmos
M$1392 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1393 r0 *1 865.09,634.52 sg13_hv_pmos
M$1393 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1394 r0 *1 865.09,635.4 sg13_hv_pmos
M$1394 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1395 r0 *1 865.09,636.28 sg13_hv_pmos
M$1395 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1396 r0 *1 865.09,637.16 sg13_hv_pmos
M$1396 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1397 r0 *1 865.09,638.04 sg13_hv_pmos
M$1397 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1398 r0 *1 865.09,638.92 sg13_hv_pmos
M$1398 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1399 r0 *1 865.09,639.8 sg13_hv_pmos
M$1399 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1400 r0 *1 865.09,640.68 sg13_hv_pmos
M$1400 IOVDD IOVDD \$626 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1401 r0 *1 865.09,641.56 sg13_hv_pmos
M$1401 \$626 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1402 r0 *1 -108.92,605.52 sg13_hv_pmos
M$1402 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1403 r0 *1 -108.92,607.3 sg13_hv_pmos
M$1403 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1404 r0 *1 -108.92,608.54 sg13_hv_pmos
M$1404 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1405 r0 *1 -108.92,610.32 sg13_hv_pmos
M$1405 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1406 r0 *1 -108.92,611.56 sg13_hv_pmos
M$1406 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1407 r0 *1 -108.92,613.34 sg13_hv_pmos
M$1407 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1408 r0 *1 -108.92,614.58 sg13_hv_pmos
M$1408 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1409 r0 *1 -108.92,616.36 sg13_hv_pmos
M$1409 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1410 r0 *1 -108.92,617.6 sg13_hv_pmos
M$1410 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1411 r0 *1 -108.92,619.38 sg13_hv_pmos
M$1411 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1412 r0 *1 -108.92,620.62 sg13_hv_pmos
M$1412 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1413 r0 *1 -108.92,622.4 sg13_hv_pmos
M$1413 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1414 r0 *1 -108.92,623.64 sg13_hv_pmos
M$1414 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1415 r0 *1 -108.92,625.42 sg13_hv_pmos
M$1415 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1416 r0 *1 -108.92,626.66 sg13_hv_pmos
M$1416 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1417 r0 *1 -108.92,628.44 sg13_hv_pmos
M$1417 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1418 r0 *1 -108.92,629.68 sg13_hv_pmos
M$1418 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1419 r0 *1 -108.92,631.46 sg13_hv_pmos
M$1419 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1420 r0 *1 -108.92,632.7 sg13_hv_pmos
M$1420 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1421 r0 *1 -108.92,634.48 sg13_hv_pmos
M$1421 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1422 r0 *1 -101.82,605.52 sg13_hv_pmos
M$1422 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1423 r0 *1 -101.82,607.3 sg13_hv_pmos
M$1423 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1424 r0 *1 -101.82,608.54 sg13_hv_pmos
M$1424 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1425 r0 *1 -101.82,610.32 sg13_hv_pmos
M$1425 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1426 r0 *1 -101.82,611.56 sg13_hv_pmos
M$1426 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1427 r0 *1 -101.82,613.34 sg13_hv_pmos
M$1427 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1428 r0 *1 -101.82,614.58 sg13_hv_pmos
M$1428 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1429 r0 *1 -101.82,616.36 sg13_hv_pmos
M$1429 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1430 r0 *1 -101.82,617.6 sg13_hv_pmos
M$1430 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1431 r0 *1 -101.82,619.38 sg13_hv_pmos
M$1431 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1432 r0 *1 -101.82,620.62 sg13_hv_pmos
M$1432 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1433 r0 *1 -101.82,622.4 sg13_hv_pmos
M$1433 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1434 r0 *1 -101.82,623.64 sg13_hv_pmos
M$1434 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1435 r0 *1 -101.82,625.42 sg13_hv_pmos
M$1435 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1436 r0 *1 -101.82,626.66 sg13_hv_pmos
M$1436 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1437 r0 *1 -101.82,628.44 sg13_hv_pmos
M$1437 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1438 r0 *1 -101.82,629.68 sg13_hv_pmos
M$1438 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1439 r0 *1 -101.82,631.46 sg13_hv_pmos
M$1439 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1440 r0 *1 -101.82,632.7 sg13_hv_pmos
M$1440 AVDD|IOVDD \$639 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1441 r0 *1 -101.82,634.48 sg13_hv_pmos
M$1441 PAD|VHI \$639 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1442 r0 *1 -108.92,705.52 sg13_hv_pmos
M$1442 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1443 r0 *1 -108.92,707.3 sg13_hv_pmos
M$1443 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1444 r0 *1 -108.92,708.54 sg13_hv_pmos
M$1444 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1445 r0 *1 -108.92,710.32 sg13_hv_pmos
M$1445 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1446 r0 *1 -108.92,711.56 sg13_hv_pmos
M$1446 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1447 r0 *1 -108.92,713.34 sg13_hv_pmos
M$1447 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1448 r0 *1 -108.92,714.58 sg13_hv_pmos
M$1448 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1449 r0 *1 -108.92,716.36 sg13_hv_pmos
M$1449 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1450 r0 *1 -108.92,717.6 sg13_hv_pmos
M$1450 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1451 r0 *1 -108.92,719.38 sg13_hv_pmos
M$1451 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1452 r0 *1 -108.92,720.62 sg13_hv_pmos
M$1452 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1453 r0 *1 -108.92,722.4 sg13_hv_pmos
M$1453 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1454 r0 *1 -108.92,723.64 sg13_hv_pmos
M$1454 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1455 r0 *1 -108.92,725.42 sg13_hv_pmos
M$1455 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1456 r0 *1 -108.92,726.66 sg13_hv_pmos
M$1456 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1457 r0 *1 -108.92,728.44 sg13_hv_pmos
M$1457 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1458 r0 *1 -108.92,729.68 sg13_hv_pmos
M$1458 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1459 r0 *1 -108.92,731.46 sg13_hv_pmos
M$1459 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1460 r0 *1 -108.92,732.7 sg13_hv_pmos
M$1460 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1461 r0 *1 -108.92,734.48 sg13_hv_pmos
M$1461 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1462 r0 *1 -101.82,705.52 sg13_hv_pmos
M$1462 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1463 r0 *1 -101.82,707.3 sg13_hv_pmos
M$1463 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1464 r0 *1 -101.82,708.54 sg13_hv_pmos
M$1464 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1465 r0 *1 -101.82,710.32 sg13_hv_pmos
M$1465 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1466 r0 *1 -101.82,711.56 sg13_hv_pmos
M$1466 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1467 r0 *1 -101.82,713.34 sg13_hv_pmos
M$1467 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1468 r0 *1 -101.82,714.58 sg13_hv_pmos
M$1468 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1469 r0 *1 -101.82,716.36 sg13_hv_pmos
M$1469 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1470 r0 *1 -101.82,717.6 sg13_hv_pmos
M$1470 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1471 r0 *1 -101.82,719.38 sg13_hv_pmos
M$1471 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1472 r0 *1 -101.82,720.62 sg13_hv_pmos
M$1472 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1473 r0 *1 -101.82,722.4 sg13_hv_pmos
M$1473 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1474 r0 *1 -101.82,723.64 sg13_hv_pmos
M$1474 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1475 r0 *1 -101.82,725.42 sg13_hv_pmos
M$1475 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1476 r0 *1 -101.82,726.66 sg13_hv_pmos
M$1476 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1477 r0 *1 -101.82,728.44 sg13_hv_pmos
M$1477 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1478 r0 *1 -101.82,729.68 sg13_hv_pmos
M$1478 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1479 r0 *1 -101.82,731.46 sg13_hv_pmos
M$1479 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1480 r0 *1 -101.82,732.7 sg13_hv_pmos
M$1480 AVDD|IOVDD \$741 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1481 r0 *1 -101.82,734.48 sg13_hv_pmos
M$1481 IN3|PAD \$741 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1482 r0 *1 881.82,714.58 sg13_hv_pmos
M$1482 IOVDD \$731 OUT3 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1483 r0 *1 881.82,716.36 sg13_hv_pmos
M$1483 OUT3 \$731 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1484 r0 *1 881.82,717.6 sg13_hv_pmos
M$1484 IOVDD \$731 OUT3 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1485 r0 *1 881.82,719.38 sg13_hv_pmos
M$1485 OUT3 \$731 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1486 r0 *1 881.82,720.62 sg13_hv_pmos
M$1486 IOVDD \$731 OUT3 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1487 r0 *1 881.82,722.4 sg13_hv_pmos
M$1487 OUT3 \$731 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1488 r0 *1 881.82,723.64 sg13_hv_pmos
M$1488 IOVDD \$731 OUT3 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1489 r0 *1 881.82,725.42 sg13_hv_pmos
M$1489 OUT3 \$731 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1490 r0 *1 888.92,714.58 sg13_hv_pmos
M$1490 IOVDD \$731 OUT3 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1491 r0 *1 888.92,716.36 sg13_hv_pmos
M$1491 OUT3 \$731 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1492 r0 *1 888.92,717.6 sg13_hv_pmos
M$1492 IOVDD \$731 OUT3 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1493 r0 *1 888.92,719.38 sg13_hv_pmos
M$1493 OUT3 \$731 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1494 r0 *1 888.92,720.62 sg13_hv_pmos
M$1494 IOVDD \$731 OUT3 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1495 r0 *1 888.92,722.4 sg13_hv_pmos
M$1495 OUT3 \$731 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1496 r0 *1 888.92,723.64 sg13_hv_pmos
M$1496 IOVDD \$731 OUT3 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1497 r0 *1 888.92,725.42 sg13_hv_pmos
M$1497 OUT3 \$731 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1498 r0 *1 808.82,717.64 sg13_hv_pmos
M$1498 \$751 \$761 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1499 r0 *1 808.82,718.47 sg13_hv_pmos
M$1499 IOVDD \$751 \$761 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1500 r0 *1 808.82,719.81 sg13_hv_pmos
M$1500 IOVDD \$761 \$766 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1501 r0 *1 808.82,721.15 sg13_hv_pmos
M$1501 \$778 \$785 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1502 r0 *1 808.82,721.98 sg13_hv_pmos
M$1502 IOVDD \$778 \$785 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1503 r0 *1 808.82,723.32 sg13_hv_pmos
M$1503 IOVDD \$785 \$731 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1504 r0 *1 -108.92,805.52 sg13_hv_pmos
M$1504 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1505 r0 *1 -108.92,807.3 sg13_hv_pmos
M$1505 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1506 r0 *1 -108.92,808.54 sg13_hv_pmos
M$1506 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1507 r0 *1 -108.92,810.32 sg13_hv_pmos
M$1507 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1508 r0 *1 -108.92,811.56 sg13_hv_pmos
M$1508 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1509 r0 *1 -108.92,813.34 sg13_hv_pmos
M$1509 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1510 r0 *1 -108.92,814.58 sg13_hv_pmos
M$1510 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1511 r0 *1 -108.92,816.36 sg13_hv_pmos
M$1511 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1512 r0 *1 -108.92,817.6 sg13_hv_pmos
M$1512 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1513 r0 *1 -108.92,819.38 sg13_hv_pmos
M$1513 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1514 r0 *1 -108.92,820.62 sg13_hv_pmos
M$1514 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1515 r0 *1 -108.92,822.4 sg13_hv_pmos
M$1515 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1516 r0 *1 -108.92,823.64 sg13_hv_pmos
M$1516 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1517 r0 *1 -108.92,825.42 sg13_hv_pmos
M$1517 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1518 r0 *1 -108.92,826.66 sg13_hv_pmos
M$1518 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1519 r0 *1 -108.92,828.44 sg13_hv_pmos
M$1519 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1520 r0 *1 -108.92,829.68 sg13_hv_pmos
M$1520 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1521 r0 *1 -108.92,831.46 sg13_hv_pmos
M$1521 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1522 r0 *1 -108.92,832.7 sg13_hv_pmos
M$1522 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1523 r0 *1 -108.92,834.48 sg13_hv_pmos
M$1523 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1524 r0 *1 -101.82,805.52 sg13_hv_pmos
M$1524 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1525 r0 *1 -101.82,807.3 sg13_hv_pmos
M$1525 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1526 r0 *1 -101.82,808.54 sg13_hv_pmos
M$1526 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1527 r0 *1 -101.82,810.32 sg13_hv_pmos
M$1527 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1528 r0 *1 -101.82,811.56 sg13_hv_pmos
M$1528 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1529 r0 *1 -101.82,813.34 sg13_hv_pmos
M$1529 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1530 r0 *1 -101.82,814.58 sg13_hv_pmos
M$1530 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1531 r0 *1 -101.82,816.36 sg13_hv_pmos
M$1531 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1532 r0 *1 -101.82,817.6 sg13_hv_pmos
M$1532 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1533 r0 *1 -101.82,819.38 sg13_hv_pmos
M$1533 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1534 r0 *1 -101.82,820.62 sg13_hv_pmos
M$1534 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1535 r0 *1 -101.82,822.4 sg13_hv_pmos
M$1535 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1536 r0 *1 -101.82,823.64 sg13_hv_pmos
M$1536 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1537 r0 *1 -101.82,825.42 sg13_hv_pmos
M$1537 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1538 r0 *1 -101.82,826.66 sg13_hv_pmos
M$1538 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1539 r0 *1 -101.82,828.44 sg13_hv_pmos
M$1539 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1540 r0 *1 -101.82,829.68 sg13_hv_pmos
M$1540 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1541 r0 *1 -101.82,831.46 sg13_hv_pmos
M$1541 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1542 r0 *1 -101.82,832.7 sg13_hv_pmos
M$1542 AVDD|IOVDD \$854 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1543 r0 *1 -101.82,834.48 sg13_hv_pmos
M$1543 IN2|PAD \$854 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1544 r0 *1 881.82,814.58 sg13_hv_pmos
M$1544 IOVDD \$844 OUT2 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1545 r0 *1 881.82,816.36 sg13_hv_pmos
M$1545 OUT2 \$844 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1546 r0 *1 881.82,817.6 sg13_hv_pmos
M$1546 IOVDD \$844 OUT2 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1547 r0 *1 881.82,819.38 sg13_hv_pmos
M$1547 OUT2 \$844 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1548 r0 *1 881.82,820.62 sg13_hv_pmos
M$1548 IOVDD \$844 OUT2 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1549 r0 *1 881.82,822.4 sg13_hv_pmos
M$1549 OUT2 \$844 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1550 r0 *1 881.82,823.64 sg13_hv_pmos
M$1550 IOVDD \$844 OUT2 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1551 r0 *1 881.82,825.42 sg13_hv_pmos
M$1551 OUT2 \$844 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1552 r0 *1 888.92,814.58 sg13_hv_pmos
M$1552 IOVDD \$844 OUT2 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1553 r0 *1 888.92,816.36 sg13_hv_pmos
M$1553 OUT2 \$844 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1554 r0 *1 888.92,817.6 sg13_hv_pmos
M$1554 IOVDD \$844 OUT2 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1555 r0 *1 888.92,819.38 sg13_hv_pmos
M$1555 OUT2 \$844 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1556 r0 *1 888.92,820.62 sg13_hv_pmos
M$1556 IOVDD \$844 OUT2 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1557 r0 *1 888.92,822.4 sg13_hv_pmos
M$1557 OUT2 \$844 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1558 r0 *1 888.92,823.64 sg13_hv_pmos
M$1558 IOVDD \$844 OUT2 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1559 r0 *1 888.92,825.42 sg13_hv_pmos
M$1559 OUT2 \$844 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1560 r0 *1 808.82,817.64 sg13_hv_pmos
M$1560 \$864 \$874 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1561 r0 *1 808.82,818.47 sg13_hv_pmos
M$1561 IOVDD \$864 \$874 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1562 r0 *1 808.82,819.81 sg13_hv_pmos
M$1562 IOVDD \$874 \$879 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1563 r0 *1 808.82,821.15 sg13_hv_pmos
M$1563 \$891 \$898 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1564 r0 *1 808.82,821.98 sg13_hv_pmos
M$1564 IOVDD \$891 \$898 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1565 r0 *1 808.82,823.32 sg13_hv_pmos
M$1565 IOVDD \$898 \$844 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1566 r0 *1 -108.92,905.52 sg13_hv_pmos
M$1566 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1567 r0 *1 -108.92,907.3 sg13_hv_pmos
M$1567 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1568 r0 *1 -108.92,908.54 sg13_hv_pmos
M$1568 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1569 r0 *1 -108.92,910.32 sg13_hv_pmos
M$1569 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1570 r0 *1 -108.92,911.56 sg13_hv_pmos
M$1570 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1571 r0 *1 -108.92,913.34 sg13_hv_pmos
M$1571 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1572 r0 *1 -108.92,914.58 sg13_hv_pmos
M$1572 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1573 r0 *1 -108.92,916.36 sg13_hv_pmos
M$1573 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1574 r0 *1 -108.92,917.6 sg13_hv_pmos
M$1574 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1575 r0 *1 -108.92,919.38 sg13_hv_pmos
M$1575 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1576 r0 *1 -108.92,920.62 sg13_hv_pmos
M$1576 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1577 r0 *1 -108.92,922.4 sg13_hv_pmos
M$1577 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1578 r0 *1 -108.92,923.64 sg13_hv_pmos
M$1578 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1579 r0 *1 -108.92,925.42 sg13_hv_pmos
M$1579 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1580 r0 *1 -108.92,926.66 sg13_hv_pmos
M$1580 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1581 r0 *1 -108.92,928.44 sg13_hv_pmos
M$1581 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1582 r0 *1 -108.92,929.68 sg13_hv_pmos
M$1582 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1583 r0 *1 -108.92,931.46 sg13_hv_pmos
M$1583 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1584 r0 *1 -108.92,932.7 sg13_hv_pmos
M$1584 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1585 r0 *1 -108.92,934.48 sg13_hv_pmos
M$1585 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1586 r0 *1 -101.82,905.52 sg13_hv_pmos
M$1586 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1587 r0 *1 -101.82,907.3 sg13_hv_pmos
M$1587 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1588 r0 *1 -101.82,908.54 sg13_hv_pmos
M$1588 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1589 r0 *1 -101.82,910.32 sg13_hv_pmos
M$1589 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1590 r0 *1 -101.82,911.56 sg13_hv_pmos
M$1590 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1591 r0 *1 -101.82,913.34 sg13_hv_pmos
M$1591 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1592 r0 *1 -101.82,914.58 sg13_hv_pmos
M$1592 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1593 r0 *1 -101.82,916.36 sg13_hv_pmos
M$1593 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1594 r0 *1 -101.82,917.6 sg13_hv_pmos
M$1594 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1595 r0 *1 -101.82,919.38 sg13_hv_pmos
M$1595 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1596 r0 *1 -101.82,920.62 sg13_hv_pmos
M$1596 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1597 r0 *1 -101.82,922.4 sg13_hv_pmos
M$1597 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1598 r0 *1 -101.82,923.64 sg13_hv_pmos
M$1598 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1599 r0 *1 -101.82,925.42 sg13_hv_pmos
M$1599 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1600 r0 *1 -101.82,926.66 sg13_hv_pmos
M$1600 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1601 r0 *1 -101.82,928.44 sg13_hv_pmos
M$1601 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1602 r0 *1 -101.82,929.68 sg13_hv_pmos
M$1602 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1603 r0 *1 -101.82,931.46 sg13_hv_pmos
M$1603 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1604 r0 *1 -101.82,932.7 sg13_hv_pmos
M$1604 AVDD|IOVDD \$967 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1605 r0 *1 -101.82,934.48 sg13_hv_pmos
M$1605 IN1|PAD \$967 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1606 r0 *1 881.82,914.58 sg13_hv_pmos
M$1606 IOVDD \$957 OUT1 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1607 r0 *1 881.82,916.36 sg13_hv_pmos
M$1607 OUT1 \$957 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1608 r0 *1 881.82,917.6 sg13_hv_pmos
M$1608 IOVDD \$957 OUT1 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1609 r0 *1 881.82,919.38 sg13_hv_pmos
M$1609 OUT1 \$957 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1610 r0 *1 881.82,920.62 sg13_hv_pmos
M$1610 IOVDD \$957 OUT1 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1611 r0 *1 881.82,922.4 sg13_hv_pmos
M$1611 OUT1 \$957 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1612 r0 *1 881.82,923.64 sg13_hv_pmos
M$1612 IOVDD \$957 OUT1 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1613 r0 *1 881.82,925.42 sg13_hv_pmos
M$1613 OUT1 \$957 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1614 r0 *1 888.92,914.58 sg13_hv_pmos
M$1614 IOVDD \$957 OUT1 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1615 r0 *1 888.92,916.36 sg13_hv_pmos
M$1615 OUT1 \$957 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1616 r0 *1 888.92,917.6 sg13_hv_pmos
M$1616 IOVDD \$957 OUT1 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1617 r0 *1 888.92,919.38 sg13_hv_pmos
M$1617 OUT1 \$957 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1618 r0 *1 888.92,920.62 sg13_hv_pmos
M$1618 IOVDD \$957 OUT1 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1619 r0 *1 888.92,922.4 sg13_hv_pmos
M$1619 OUT1 \$957 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1620 r0 *1 888.92,923.64 sg13_hv_pmos
M$1620 IOVDD \$957 OUT1 IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1621 r0 *1 888.92,925.42 sg13_hv_pmos
M$1621 OUT1 \$957 IOVDD IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1622 r0 *1 808.82,917.64 sg13_hv_pmos
M$1622 \$977 \$987 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1623 r0 *1 808.82,918.47 sg13_hv_pmos
M$1623 IOVDD \$977 \$987 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1624 r0 *1 808.82,919.81 sg13_hv_pmos
M$1624 IOVDD \$987 \$992 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1625 r0 *1 808.82,921.15 sg13_hv_pmos
M$1625 \$1004 \$1011 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1626 r0 *1 808.82,921.98 sg13_hv_pmos
M$1626 IOVDD \$1004 \$1011 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1627 r0 *1 808.82,923.32 sg13_hv_pmos
M$1627 IOVDD \$1011 \$957 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1628 r0 *1 441.765,976.055 sg13_hv_pmos
M$1628 VDD \$1070 \$1067 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1629 r0 *1 541.765,976.055 sg13_hv_pmos
M$1629 VDD \$1071 \$1068 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1630 r0 *1 641.765,976.055 sg13_hv_pmos
M$1630 VDD \$1072 \$1069 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1631 r0 *1 18.44,1045.09 sg13_hv_pmos
M$1631 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1632 r0 *1 19.32,1045.09 sg13_hv_pmos
M$1632 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1633 r0 *1 20.2,1045.09 sg13_hv_pmos
M$1633 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1634 r0 *1 21.08,1045.09 sg13_hv_pmos
M$1634 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1635 r0 *1 21.96,1045.09 sg13_hv_pmos
M$1635 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1636 r0 *1 22.84,1045.09 sg13_hv_pmos
M$1636 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1637 r0 *1 23.72,1045.09 sg13_hv_pmos
M$1637 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1638 r0 *1 24.6,1045.09 sg13_hv_pmos
M$1638 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1639 r0 *1 25.48,1045.09 sg13_hv_pmos
M$1639 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1640 r0 *1 26.36,1045.09 sg13_hv_pmos
M$1640 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1641 r0 *1 27.24,1045.09 sg13_hv_pmos
M$1641 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1642 r0 *1 28.12,1045.09 sg13_hv_pmos
M$1642 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1643 r0 *1 29,1045.09 sg13_hv_pmos
M$1643 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1644 r0 *1 29.88,1045.09 sg13_hv_pmos
M$1644 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1645 r0 *1 30.76,1045.09 sg13_hv_pmos
M$1645 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1646 r0 *1 31.64,1045.09 sg13_hv_pmos
M$1646 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1647 r0 *1 32.52,1045.09 sg13_hv_pmos
M$1647 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1648 r0 *1 33.4,1045.09 sg13_hv_pmos
M$1648 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1649 r0 *1 34.28,1045.09 sg13_hv_pmos
M$1649 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1650 r0 *1 35.16,1045.09 sg13_hv_pmos
M$1650 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1651 r0 *1 36.04,1045.09 sg13_hv_pmos
M$1651 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1652 r0 *1 36.92,1045.09 sg13_hv_pmos
M$1652 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1653 r0 *1 37.8,1045.09 sg13_hv_pmos
M$1653 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1654 r0 *1 38.68,1045.09 sg13_hv_pmos
M$1654 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1655 r0 *1 39.56,1045.09 sg13_hv_pmos
M$1655 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1656 r0 *1 40.44,1045.09 sg13_hv_pmos
M$1656 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1657 r0 *1 41.32,1045.09 sg13_hv_pmos
M$1657 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1658 r0 *1 42.2,1045.09 sg13_hv_pmos
M$1658 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1659 r0 *1 43.08,1045.09 sg13_hv_pmos
M$1659 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1660 r0 *1 43.96,1045.09 sg13_hv_pmos
M$1660 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1661 r0 *1 44.84,1045.09 sg13_hv_pmos
M$1661 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1662 r0 *1 45.72,1045.09 sg13_hv_pmos
M$1662 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1663 r0 *1 46.6,1045.09 sg13_hv_pmos
M$1663 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1664 r0 *1 47.48,1045.09 sg13_hv_pmos
M$1664 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1665 r0 *1 48.36,1045.09 sg13_hv_pmos
M$1665 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1666 r0 *1 49.24,1045.09 sg13_hv_pmos
M$1666 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1667 r0 *1 50.12,1045.09 sg13_hv_pmos
M$1667 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1668 r0 *1 51,1045.09 sg13_hv_pmos
M$1668 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1669 r0 *1 51.88,1045.09 sg13_hv_pmos
M$1669 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1670 r0 *1 52.76,1045.09 sg13_hv_pmos
M$1670 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1671 r0 *1 53.64,1045.09 sg13_hv_pmos
M$1671 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1672 r0 *1 54.52,1045.09 sg13_hv_pmos
M$1672 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1673 r0 *1 55.4,1045.09 sg13_hv_pmos
M$1673 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1674 r0 *1 56.28,1045.09 sg13_hv_pmos
M$1674 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1675 r0 *1 57.16,1045.09 sg13_hv_pmos
M$1675 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1676 r0 *1 58.04,1045.09 sg13_hv_pmos
M$1676 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1677 r0 *1 58.92,1045.09 sg13_hv_pmos
M$1677 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1678 r0 *1 59.8,1045.09 sg13_hv_pmos
M$1678 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1679 r0 *1 60.68,1045.09 sg13_hv_pmos
M$1679 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1680 r0 *1 61.56,1045.09 sg13_hv_pmos
M$1680 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1681 r0 *1 318.44,1045.09 sg13_hv_pmos
M$1681 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1682 r0 *1 319.32,1045.09 sg13_hv_pmos
M$1682 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1683 r0 *1 320.2,1045.09 sg13_hv_pmos
M$1683 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1684 r0 *1 321.08,1045.09 sg13_hv_pmos
M$1684 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1685 r0 *1 321.96,1045.09 sg13_hv_pmos
M$1685 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1686 r0 *1 322.84,1045.09 sg13_hv_pmos
M$1686 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1687 r0 *1 323.72,1045.09 sg13_hv_pmos
M$1687 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1688 r0 *1 324.6,1045.09 sg13_hv_pmos
M$1688 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1689 r0 *1 325.48,1045.09 sg13_hv_pmos
M$1689 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1690 r0 *1 326.36,1045.09 sg13_hv_pmos
M$1690 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1691 r0 *1 327.24,1045.09 sg13_hv_pmos
M$1691 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1692 r0 *1 328.12,1045.09 sg13_hv_pmos
M$1692 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1693 r0 *1 329,1045.09 sg13_hv_pmos
M$1693 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1694 r0 *1 329.88,1045.09 sg13_hv_pmos
M$1694 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1695 r0 *1 330.76,1045.09 sg13_hv_pmos
M$1695 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1696 r0 *1 331.64,1045.09 sg13_hv_pmos
M$1696 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1697 r0 *1 332.52,1045.09 sg13_hv_pmos
M$1697 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1698 r0 *1 333.4,1045.09 sg13_hv_pmos
M$1698 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1699 r0 *1 334.28,1045.09 sg13_hv_pmos
M$1699 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1700 r0 *1 335.16,1045.09 sg13_hv_pmos
M$1700 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1701 r0 *1 336.04,1045.09 sg13_hv_pmos
M$1701 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1702 r0 *1 336.92,1045.09 sg13_hv_pmos
M$1702 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1703 r0 *1 337.8,1045.09 sg13_hv_pmos
M$1703 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1704 r0 *1 338.68,1045.09 sg13_hv_pmos
M$1704 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1705 r0 *1 339.56,1045.09 sg13_hv_pmos
M$1705 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1706 r0 *1 340.44,1045.09 sg13_hv_pmos
M$1706 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1707 r0 *1 341.32,1045.09 sg13_hv_pmos
M$1707 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1708 r0 *1 342.2,1045.09 sg13_hv_pmos
M$1708 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1709 r0 *1 343.08,1045.09 sg13_hv_pmos
M$1709 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1710 r0 *1 343.96,1045.09 sg13_hv_pmos
M$1710 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1711 r0 *1 344.84,1045.09 sg13_hv_pmos
M$1711 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1712 r0 *1 345.72,1045.09 sg13_hv_pmos
M$1712 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1713 r0 *1 346.6,1045.09 sg13_hv_pmos
M$1713 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1714 r0 *1 347.48,1045.09 sg13_hv_pmos
M$1714 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1715 r0 *1 348.36,1045.09 sg13_hv_pmos
M$1715 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1716 r0 *1 349.24,1045.09 sg13_hv_pmos
M$1716 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1717 r0 *1 350.12,1045.09 sg13_hv_pmos
M$1717 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1718 r0 *1 351,1045.09 sg13_hv_pmos
M$1718 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1719 r0 *1 351.88,1045.09 sg13_hv_pmos
M$1719 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1720 r0 *1 352.76,1045.09 sg13_hv_pmos
M$1720 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1721 r0 *1 353.64,1045.09 sg13_hv_pmos
M$1721 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1722 r0 *1 354.52,1045.09 sg13_hv_pmos
M$1722 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1723 r0 *1 355.4,1045.09 sg13_hv_pmos
M$1723 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1724 r0 *1 356.28,1045.09 sg13_hv_pmos
M$1724 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1725 r0 *1 357.16,1045.09 sg13_hv_pmos
M$1725 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1726 r0 *1 358.04,1045.09 sg13_hv_pmos
M$1726 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1727 r0 *1 358.92,1045.09 sg13_hv_pmos
M$1727 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1728 r0 *1 359.8,1045.09 sg13_hv_pmos
M$1728 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1729 r0 *1 360.68,1045.09 sg13_hv_pmos
M$1729 IOVDD IOVDD \$1144 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1730 r0 *1 361.56,1045.09 sg13_hv_pmos
M$1730 \$1144 IOVDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1731 r0 *1 718.44,1045.09 sg13_hv_pmos
M$1731 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1732 r0 *1 719.32,1045.09 sg13_hv_pmos
M$1732 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1733 r0 *1 720.2,1045.09 sg13_hv_pmos
M$1733 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1734 r0 *1 721.08,1045.09 sg13_hv_pmos
M$1734 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1735 r0 *1 721.96,1045.09 sg13_hv_pmos
M$1735 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1736 r0 *1 722.84,1045.09 sg13_hv_pmos
M$1736 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1737 r0 *1 723.72,1045.09 sg13_hv_pmos
M$1737 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1738 r0 *1 724.6,1045.09 sg13_hv_pmos
M$1738 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1739 r0 *1 725.48,1045.09 sg13_hv_pmos
M$1739 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1740 r0 *1 726.36,1045.09 sg13_hv_pmos
M$1740 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1741 r0 *1 727.24,1045.09 sg13_hv_pmos
M$1741 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1742 r0 *1 728.12,1045.09 sg13_hv_pmos
M$1742 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1743 r0 *1 729,1045.09 sg13_hv_pmos
M$1743 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1744 r0 *1 729.88,1045.09 sg13_hv_pmos
M$1744 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1745 r0 *1 730.76,1045.09 sg13_hv_pmos
M$1745 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1746 r0 *1 731.64,1045.09 sg13_hv_pmos
M$1746 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1747 r0 *1 732.52,1045.09 sg13_hv_pmos
M$1747 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1748 r0 *1 733.4,1045.09 sg13_hv_pmos
M$1748 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1749 r0 *1 734.28,1045.09 sg13_hv_pmos
M$1749 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1750 r0 *1 735.16,1045.09 sg13_hv_pmos
M$1750 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1751 r0 *1 736.04,1045.09 sg13_hv_pmos
M$1751 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1752 r0 *1 736.92,1045.09 sg13_hv_pmos
M$1752 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1753 r0 *1 737.8,1045.09 sg13_hv_pmos
M$1753 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1754 r0 *1 738.68,1045.09 sg13_hv_pmos
M$1754 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1755 r0 *1 739.56,1045.09 sg13_hv_pmos
M$1755 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1756 r0 *1 740.44,1045.09 sg13_hv_pmos
M$1756 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1757 r0 *1 741.32,1045.09 sg13_hv_pmos
M$1757 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1758 r0 *1 742.2,1045.09 sg13_hv_pmos
M$1758 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1759 r0 *1 743.08,1045.09 sg13_hv_pmos
M$1759 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1760 r0 *1 743.96,1045.09 sg13_hv_pmos
M$1760 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1761 r0 *1 744.84,1045.09 sg13_hv_pmos
M$1761 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1762 r0 *1 745.72,1045.09 sg13_hv_pmos
M$1762 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1763 r0 *1 746.6,1045.09 sg13_hv_pmos
M$1763 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1764 r0 *1 747.48,1045.09 sg13_hv_pmos
M$1764 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1765 r0 *1 748.36,1045.09 sg13_hv_pmos
M$1765 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1766 r0 *1 749.24,1045.09 sg13_hv_pmos
M$1766 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1767 r0 *1 750.12,1045.09 sg13_hv_pmos
M$1767 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1768 r0 *1 751,1045.09 sg13_hv_pmos
M$1768 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1769 r0 *1 751.88,1045.09 sg13_hv_pmos
M$1769 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1770 r0 *1 752.76,1045.09 sg13_hv_pmos
M$1770 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1771 r0 *1 753.64,1045.09 sg13_hv_pmos
M$1771 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1772 r0 *1 754.52,1045.09 sg13_hv_pmos
M$1772 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1773 r0 *1 755.4,1045.09 sg13_hv_pmos
M$1773 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1774 r0 *1 756.28,1045.09 sg13_hv_pmos
M$1774 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1775 r0 *1 757.16,1045.09 sg13_hv_pmos
M$1775 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1776 r0 *1 758.04,1045.09 sg13_hv_pmos
M$1776 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1777 r0 *1 758.92,1045.09 sg13_hv_pmos
M$1777 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1778 r0 *1 759.8,1045.09 sg13_hv_pmos
M$1778 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1779 r0 *1 760.68,1045.09 sg13_hv_pmos
M$1779 IOVDD VDD \$1145 IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1780 r0 *1 761.56,1045.09 sg13_hv_pmos
M$1780 \$1145 VDD IOVDD IOVDD sg13_hv_pmos W=6.999999999999998
+ L=0.4999999999999999
* device instance $1781 r0 *1 125.52,1061.82 sg13_hv_pmos
M$1781 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1782 r0 *1 127.3,1061.82 sg13_hv_pmos
M$1782 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1783 r0 *1 128.54,1061.82 sg13_hv_pmos
M$1783 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1784 r0 *1 130.32,1061.82 sg13_hv_pmos
M$1784 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1785 r0 *1 131.56,1061.82 sg13_hv_pmos
M$1785 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1786 r0 *1 133.34,1061.82 sg13_hv_pmos
M$1786 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1787 r0 *1 134.58,1061.82 sg13_hv_pmos
M$1787 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1788 r0 *1 136.36,1061.82 sg13_hv_pmos
M$1788 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1789 r0 *1 137.6,1061.82 sg13_hv_pmos
M$1789 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1790 r0 *1 139.38,1061.82 sg13_hv_pmos
M$1790 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1791 r0 *1 140.62,1061.82 sg13_hv_pmos
M$1791 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1792 r0 *1 142.4,1061.82 sg13_hv_pmos
M$1792 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1793 r0 *1 143.64,1061.82 sg13_hv_pmos
M$1793 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1794 r0 *1 145.42,1061.82 sg13_hv_pmos
M$1794 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1795 r0 *1 146.66,1061.82 sg13_hv_pmos
M$1795 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1796 r0 *1 148.44,1061.82 sg13_hv_pmos
M$1796 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1797 r0 *1 149.68,1061.82 sg13_hv_pmos
M$1797 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1798 r0 *1 151.46,1061.82 sg13_hv_pmos
M$1798 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1799 r0 *1 152.7,1061.82 sg13_hv_pmos
M$1799 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1800 r0 *1 154.48,1061.82 sg13_hv_pmos
M$1800 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1801 r0 *1 125.52,1068.92 sg13_hv_pmos
M$1801 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1802 r0 *1 127.3,1068.92 sg13_hv_pmos
M$1802 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1803 r0 *1 128.54,1068.92 sg13_hv_pmos
M$1803 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1804 r0 *1 130.32,1068.92 sg13_hv_pmos
M$1804 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1805 r0 *1 131.56,1068.92 sg13_hv_pmos
M$1805 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1806 r0 *1 133.34,1068.92 sg13_hv_pmos
M$1806 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1807 r0 *1 134.58,1068.92 sg13_hv_pmos
M$1807 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1808 r0 *1 136.36,1068.92 sg13_hv_pmos
M$1808 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1809 r0 *1 137.6,1068.92 sg13_hv_pmos
M$1809 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1810 r0 *1 139.38,1068.92 sg13_hv_pmos
M$1810 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1811 r0 *1 140.62,1068.92 sg13_hv_pmos
M$1811 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1812 r0 *1 142.4,1068.92 sg13_hv_pmos
M$1812 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1813 r0 *1 143.64,1068.92 sg13_hv_pmos
M$1813 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1814 r0 *1 145.42,1068.92 sg13_hv_pmos
M$1814 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1815 r0 *1 146.66,1068.92 sg13_hv_pmos
M$1815 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1816 r0 *1 148.44,1068.92 sg13_hv_pmos
M$1816 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1817 r0 *1 149.68,1068.92 sg13_hv_pmos
M$1817 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1818 r0 *1 151.46,1068.92 sg13_hv_pmos
M$1818 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1819 r0 *1 152.7,1068.92 sg13_hv_pmos
M$1819 AVDD|IOVDD \$1160 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1820 r0 *1 154.48,1068.92 sg13_hv_pmos
M$1820 PAD|VREF \$1160 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1821 r0 *1 225.52,1061.82 sg13_hv_pmos
M$1821 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1822 r0 *1 227.3,1061.82 sg13_hv_pmos
M$1822 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1823 r0 *1 228.54,1061.82 sg13_hv_pmos
M$1823 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1824 r0 *1 230.32,1061.82 sg13_hv_pmos
M$1824 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1825 r0 *1 231.56,1061.82 sg13_hv_pmos
M$1825 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1826 r0 *1 233.34,1061.82 sg13_hv_pmos
M$1826 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1827 r0 *1 234.58,1061.82 sg13_hv_pmos
M$1827 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1828 r0 *1 236.36,1061.82 sg13_hv_pmos
M$1828 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1829 r0 *1 237.6,1061.82 sg13_hv_pmos
M$1829 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1830 r0 *1 239.38,1061.82 sg13_hv_pmos
M$1830 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1831 r0 *1 240.62,1061.82 sg13_hv_pmos
M$1831 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1832 r0 *1 242.4,1061.82 sg13_hv_pmos
M$1832 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1833 r0 *1 243.64,1061.82 sg13_hv_pmos
M$1833 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1834 r0 *1 245.42,1061.82 sg13_hv_pmos
M$1834 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1835 r0 *1 246.66,1061.82 sg13_hv_pmos
M$1835 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1836 r0 *1 248.44,1061.82 sg13_hv_pmos
M$1836 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1837 r0 *1 249.68,1061.82 sg13_hv_pmos
M$1837 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1838 r0 *1 251.46,1061.82 sg13_hv_pmos
M$1838 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1839 r0 *1 252.7,1061.82 sg13_hv_pmos
M$1839 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1840 r0 *1 254.48,1061.82 sg13_hv_pmos
M$1840 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1841 r0 *1 225.52,1068.92 sg13_hv_pmos
M$1841 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1842 r0 *1 227.3,1068.92 sg13_hv_pmos
M$1842 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1843 r0 *1 228.54,1068.92 sg13_hv_pmos
M$1843 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1844 r0 *1 230.32,1068.92 sg13_hv_pmos
M$1844 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1845 r0 *1 231.56,1068.92 sg13_hv_pmos
M$1845 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1846 r0 *1 233.34,1068.92 sg13_hv_pmos
M$1846 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1847 r0 *1 234.58,1068.92 sg13_hv_pmos
M$1847 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1848 r0 *1 236.36,1068.92 sg13_hv_pmos
M$1848 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1849 r0 *1 237.6,1068.92 sg13_hv_pmos
M$1849 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1850 r0 *1 239.38,1068.92 sg13_hv_pmos
M$1850 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1851 r0 *1 240.62,1068.92 sg13_hv_pmos
M$1851 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1852 r0 *1 242.4,1068.92 sg13_hv_pmos
M$1852 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1853 r0 *1 243.64,1068.92 sg13_hv_pmos
M$1853 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1854 r0 *1 245.42,1068.92 sg13_hv_pmos
M$1854 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1855 r0 *1 246.66,1068.92 sg13_hv_pmos
M$1855 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1856 r0 *1 248.44,1068.92 sg13_hv_pmos
M$1856 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1857 r0 *1 249.68,1068.92 sg13_hv_pmos
M$1857 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1858 r0 *1 251.46,1068.92 sg13_hv_pmos
M$1858 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1859 r0 *1 252.7,1068.92 sg13_hv_pmos
M$1859 AVDD|IOVDD \$1161 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1860 r0 *1 254.48,1068.92 sg13_hv_pmos
M$1860 PAD|VLDO \$1161 AVDD|IOVDD AVDD|IOVDD sg13_hv_pmos W=6.659999999999998
+ L=0.5999999999999999
* device instance $1861 r0 *1 879.21,583.22 rfnmoshv
1861$1861 IOVSS|VSS IOVDD \$626 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $1862 r0 *1 879.21,584.1 rfnmoshv
1862$1862 \$626 IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $1863 r0 *1 879.21,584.98 rfnmoshv
1863$1863 IOVSS|VSS IOVDD \$626 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $1864 r0 *1 879.21,585.86 rfnmoshv
1864$1864 \$626 IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $1865 r0 *1 879.21,586.74 rfnmoshv
1865$1865 IOVSS|VSS IOVDD \$626 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $1866 r0 *1 879.21,587.62 rfnmoshv
1866$1866 \$626 IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $1867 r0 *1 879.21,593 rfnmoshv
1867$1867 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $1868 r0 *1 879.21,602.88 rfnmoshv
1868$1868 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $1869 r0 *1 879.21,612.76 rfnmoshv
1869$1869 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $1870 r0 *1 879.21,622.64 rfnmoshv
1870$1870 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $1871 r0 *1 879.21,632.52 rfnmoshv
1871$1871 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $1872 r0 *1 879.21,642.4 rfnmoshv
1872$1872 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $1873 r0 *1 879.21,652.28 rfnmoshv
1873$1873 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $1874 r0 *1 888.46,583.22 rfnmoshv
1874$1874 IOVSS|VSS IOVDD \$626 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $1875 r0 *1 888.46,584.1 rfnmoshv
1875$1875 \$626 IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $1876 r0 *1 888.46,584.98 rfnmoshv
1876$1876 IOVSS|VSS IOVDD \$626 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $1877 r0 *1 888.46,585.86 rfnmoshv
1877$1877 \$626 IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $1878 r0 *1 888.46,586.74 rfnmoshv
1878$1878 IOVSS|VSS IOVDD \$626 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $1879 r0 *1 888.46,587.62 rfnmoshv
1879$1879 \$626 IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $1880 r0 *1 888.46,593 rfnmoshv
1880$1880 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $1881 r0 *1 888.46,602.88 rfnmoshv
1881$1881 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $1882 r0 *1 888.46,612.76 rfnmoshv
1882$1882 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $1883 r0 *1 888.46,622.64 rfnmoshv
1883$1883 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $1884 r0 *1 888.46,632.52 rfnmoshv
1884$1884 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $1885 r0 *1 888.46,642.4 rfnmoshv
1885$1885 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $1886 r0 *1 888.46,652.28 rfnmoshv
1886$1886 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $1887 r0 *1 934.53,588.155 rfnmoshv
1887$1887 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1888 r0 *1 934.53,589.935 rfnmoshv
1888$1888 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1889 r0 *1 934.53,591.175 rfnmoshv
1889$1889 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1890 r0 *1 934.53,592.955 rfnmoshv
1890$1890 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1891 r0 *1 934.53,594.195 rfnmoshv
1891$1891 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1892 r0 *1 934.53,595.975 rfnmoshv
1892$1892 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1893 r0 *1 934.53,597.215 rfnmoshv
1893$1893 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1894 r0 *1 934.53,598.995 rfnmoshv
1894$1894 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1895 r0 *1 934.53,600.235 rfnmoshv
1895$1895 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1896 r0 *1 934.53,602.015 rfnmoshv
1896$1896 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1897 r0 *1 934.53,603.255 rfnmoshv
1897$1897 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1898 r0 *1 934.53,605.035 rfnmoshv
1898$1898 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1899 r0 *1 934.53,606.275 rfnmoshv
1899$1899 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1900 r0 *1 934.53,608.055 rfnmoshv
1900$1900 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1901 r0 *1 934.53,609.295 rfnmoshv
1901$1901 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1902 r0 *1 934.53,611.075 rfnmoshv
1902$1902 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1903 r0 *1 934.53,612.315 rfnmoshv
1903$1903 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1904 r0 *1 934.53,614.095 rfnmoshv
1904$1904 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1905 r0 *1 934.53,615.335 rfnmoshv
1905$1905 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1906 r0 *1 934.53,617.115 rfnmoshv
1906$1906 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1907 r0 *1 934.53,618.355 rfnmoshv
1907$1907 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1908 r0 *1 934.53,620.135 rfnmoshv
1908$1908 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1909 r0 *1 934.53,621.375 rfnmoshv
1909$1909 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1910 r0 *1 934.53,623.155 rfnmoshv
1910$1910 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1911 r0 *1 934.53,624.395 rfnmoshv
1911$1911 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1912 r0 *1 934.53,626.175 rfnmoshv
1912$1912 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1913 r0 *1 934.53,627.415 rfnmoshv
1913$1913 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1914 r0 *1 934.53,629.195 rfnmoshv
1914$1914 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1915 r0 *1 934.53,630.435 rfnmoshv
1915$1915 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1916 r0 *1 934.53,632.215 rfnmoshv
1916$1916 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1917 r0 *1 934.53,633.455 rfnmoshv
1917$1917 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1918 r0 *1 934.53,635.235 rfnmoshv
1918$1918 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1919 r0 *1 934.53,636.475 rfnmoshv
1919$1919 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1920 r0 *1 934.53,638.255 rfnmoshv
1920$1920 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1921 r0 *1 934.53,639.495 rfnmoshv
1921$1921 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1922 r0 *1 934.53,641.275 rfnmoshv
1922$1922 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1923 r0 *1 934.53,642.515 rfnmoshv
1923$1923 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1924 r0 *1 934.53,644.295 rfnmoshv
1924$1924 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1925 r0 *1 934.53,645.535 rfnmoshv
1925$1925 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1926 r0 *1 934.53,647.315 rfnmoshv
1926$1926 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1927 r0 *1 934.53,648.555 rfnmoshv
1927$1927 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1928 r0 *1 934.53,650.335 rfnmoshv
1928$1928 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1929 r0 *1 934.53,651.575 rfnmoshv
1929$1929 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1930 r0 *1 939.37,588.155 rfnmoshv
1930$1930 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1931 r0 *1 939.37,589.935 rfnmoshv
1931$1931 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1932 r0 *1 939.37,591.175 rfnmoshv
1932$1932 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1933 r0 *1 939.37,592.955 rfnmoshv
1933$1933 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1934 r0 *1 939.37,594.195 rfnmoshv
1934$1934 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1935 r0 *1 939.37,595.975 rfnmoshv
1935$1935 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1936 r0 *1 939.37,597.215 rfnmoshv
1936$1936 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1937 r0 *1 939.37,598.995 rfnmoshv
1937$1937 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1938 r0 *1 939.37,600.235 rfnmoshv
1938$1938 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1939 r0 *1 939.37,602.015 rfnmoshv
1939$1939 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1940 r0 *1 939.37,603.255 rfnmoshv
1940$1940 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1941 r0 *1 939.37,605.035 rfnmoshv
1941$1941 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1942 r0 *1 939.37,606.275 rfnmoshv
1942$1942 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1943 r0 *1 939.37,608.055 rfnmoshv
1943$1943 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1944 r0 *1 939.37,609.295 rfnmoshv
1944$1944 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1945 r0 *1 939.37,611.075 rfnmoshv
1945$1945 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1946 r0 *1 939.37,612.315 rfnmoshv
1946$1946 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1947 r0 *1 939.37,614.095 rfnmoshv
1947$1947 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1948 r0 *1 939.37,615.335 rfnmoshv
1948$1948 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1949 r0 *1 939.37,617.115 rfnmoshv
1949$1949 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1950 r0 *1 939.37,618.355 rfnmoshv
1950$1950 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1951 r0 *1 939.37,620.135 rfnmoshv
1951$1951 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1952 r0 *1 939.37,621.375 rfnmoshv
1952$1952 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1953 r0 *1 939.37,623.155 rfnmoshv
1953$1953 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1954 r0 *1 939.37,624.395 rfnmoshv
1954$1954 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1955 r0 *1 939.37,626.175 rfnmoshv
1955$1955 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1956 r0 *1 939.37,627.415 rfnmoshv
1956$1956 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1957 r0 *1 939.37,629.195 rfnmoshv
1957$1957 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1958 r0 *1 939.37,630.435 rfnmoshv
1958$1958 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1959 r0 *1 939.37,632.215 rfnmoshv
1959$1959 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1960 r0 *1 939.37,633.455 rfnmoshv
1960$1960 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1961 r0 *1 939.37,635.235 rfnmoshv
1961$1961 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1962 r0 *1 939.37,636.475 rfnmoshv
1962$1962 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1963 r0 *1 939.37,638.255 rfnmoshv
1963$1963 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1964 r0 *1 939.37,639.495 rfnmoshv
1964$1964 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1965 r0 *1 939.37,641.275 rfnmoshv
1965$1965 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1966 r0 *1 939.37,642.515 rfnmoshv
1966$1966 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1967 r0 *1 939.37,644.295 rfnmoshv
1967$1967 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1968 r0 *1 939.37,645.535 rfnmoshv
1968$1968 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1969 r0 *1 939.37,647.315 rfnmoshv
1969$1969 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1970 r0 *1 939.37,648.555 rfnmoshv
1970$1970 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1971 r0 *1 939.37,650.335 rfnmoshv
1971$1971 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1972 r0 *1 939.37,651.575 rfnmoshv
1972$1972 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1973 r0 *1 944.21,588.155 rfnmoshv
1973$1973 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1974 r0 *1 944.21,589.935 rfnmoshv
1974$1974 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1975 r0 *1 944.21,591.175 rfnmoshv
1975$1975 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1976 r0 *1 944.21,592.955 rfnmoshv
1976$1976 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1977 r0 *1 944.21,594.195 rfnmoshv
1977$1977 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1978 r0 *1 944.21,595.975 rfnmoshv
1978$1978 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1979 r0 *1 944.21,597.215 rfnmoshv
1979$1979 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1980 r0 *1 944.21,598.995 rfnmoshv
1980$1980 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1981 r0 *1 944.21,600.235 rfnmoshv
1981$1981 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1982 r0 *1 944.21,602.015 rfnmoshv
1982$1982 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1983 r0 *1 944.21,603.255 rfnmoshv
1983$1983 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1984 r0 *1 944.21,605.035 rfnmoshv
1984$1984 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1985 r0 *1 944.21,606.275 rfnmoshv
1985$1985 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1986 r0 *1 944.21,608.055 rfnmoshv
1986$1986 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1987 r0 *1 944.21,609.295 rfnmoshv
1987$1987 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1988 r0 *1 944.21,611.075 rfnmoshv
1988$1988 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1989 r0 *1 944.21,612.315 rfnmoshv
1989$1989 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1990 r0 *1 944.21,614.095 rfnmoshv
1990$1990 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1991 r0 *1 944.21,615.335 rfnmoshv
1991$1991 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1992 r0 *1 944.21,617.115 rfnmoshv
1992$1992 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1993 r0 *1 944.21,618.355 rfnmoshv
1993$1993 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1994 r0 *1 944.21,620.135 rfnmoshv
1994$1994 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1995 r0 *1 944.21,621.375 rfnmoshv
1995$1995 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1996 r0 *1 944.21,623.155 rfnmoshv
1996$1996 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1997 r0 *1 944.21,624.395 rfnmoshv
1997$1997 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1998 r0 *1 944.21,626.175 rfnmoshv
1998$1998 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $1999 r0 *1 944.21,627.415 rfnmoshv
1999$1999 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2000 r0 *1 944.21,629.195 rfnmoshv
2000$2000 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2001 r0 *1 944.21,630.435 rfnmoshv
2001$2001 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2002 r0 *1 944.21,632.215 rfnmoshv
2002$2002 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2003 r0 *1 944.21,633.455 rfnmoshv
2003$2003 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2004 r0 *1 944.21,635.235 rfnmoshv
2004$2004 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2005 r0 *1 944.21,636.475 rfnmoshv
2005$2005 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2006 r0 *1 944.21,638.255 rfnmoshv
2006$2006 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2007 r0 *1 944.21,639.495 rfnmoshv
2007$2007 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2008 r0 *1 944.21,641.275 rfnmoshv
2008$2008 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2009 r0 *1 944.21,642.515 rfnmoshv
2009$2009 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2010 r0 *1 944.21,644.295 rfnmoshv
2010$2010 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2011 r0 *1 944.21,645.535 rfnmoshv
2011$2011 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2012 r0 *1 944.21,647.315 rfnmoshv
2012$2012 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2013 r0 *1 944.21,648.555 rfnmoshv
2013$2013 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2014 r0 *1 944.21,650.335 rfnmoshv
2014$2014 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2015 r0 *1 944.21,651.575 rfnmoshv
2015$2015 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2016 r0 *1 949.05,588.155 rfnmoshv
2016$2016 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2017 r0 *1 949.05,589.935 rfnmoshv
2017$2017 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2018 r0 *1 949.05,591.175 rfnmoshv
2018$2018 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2019 r0 *1 949.05,592.955 rfnmoshv
2019$2019 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2020 r0 *1 949.05,594.195 rfnmoshv
2020$2020 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2021 r0 *1 949.05,595.975 rfnmoshv
2021$2021 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2022 r0 *1 949.05,597.215 rfnmoshv
2022$2022 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2023 r0 *1 949.05,598.995 rfnmoshv
2023$2023 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2024 r0 *1 949.05,600.235 rfnmoshv
2024$2024 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2025 r0 *1 949.05,602.015 rfnmoshv
2025$2025 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2026 r0 *1 949.05,603.255 rfnmoshv
2026$2026 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2027 r0 *1 949.05,605.035 rfnmoshv
2027$2027 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2028 r0 *1 949.05,606.275 rfnmoshv
2028$2028 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2029 r0 *1 949.05,608.055 rfnmoshv
2029$2029 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2030 r0 *1 949.05,609.295 rfnmoshv
2030$2030 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2031 r0 *1 949.05,611.075 rfnmoshv
2031$2031 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2032 r0 *1 949.05,612.315 rfnmoshv
2032$2032 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2033 r0 *1 949.05,614.095 rfnmoshv
2033$2033 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2034 r0 *1 949.05,615.335 rfnmoshv
2034$2034 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2035 r0 *1 949.05,617.115 rfnmoshv
2035$2035 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2036 r0 *1 949.05,618.355 rfnmoshv
2036$2036 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2037 r0 *1 949.05,620.135 rfnmoshv
2037$2037 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2038 r0 *1 949.05,621.375 rfnmoshv
2038$2038 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2039 r0 *1 949.05,623.155 rfnmoshv
2039$2039 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2040 r0 *1 949.05,624.395 rfnmoshv
2040$2040 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2041 r0 *1 949.05,626.175 rfnmoshv
2041$2041 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2042 r0 *1 949.05,627.415 rfnmoshv
2042$2042 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2043 r0 *1 949.05,629.195 rfnmoshv
2043$2043 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2044 r0 *1 949.05,630.435 rfnmoshv
2044$2044 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2045 r0 *1 949.05,632.215 rfnmoshv
2045$2045 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2046 r0 *1 949.05,633.455 rfnmoshv
2046$2046 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2047 r0 *1 949.05,635.235 rfnmoshv
2047$2047 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2048 r0 *1 949.05,636.475 rfnmoshv
2048$2048 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2049 r0 *1 949.05,638.255 rfnmoshv
2049$2049 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2050 r0 *1 949.05,639.495 rfnmoshv
2050$2050 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2051 r0 *1 949.05,641.275 rfnmoshv
2051$2051 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2052 r0 *1 949.05,642.515 rfnmoshv
2052$2052 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2053 r0 *1 949.05,644.295 rfnmoshv
2053$2053 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2054 r0 *1 949.05,645.535 rfnmoshv
2054$2054 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2055 r0 *1 949.05,647.315 rfnmoshv
2055$2055 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2056 r0 *1 949.05,648.555 rfnmoshv
2056$2056 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2057 r0 *1 949.05,650.335 rfnmoshv
2057$2057 IOVDD \$626 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2058 r0 *1 949.05,651.575 rfnmoshv
2058$2058 IOVSS|VSS \$626 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2059 r0 *1 3.22,1059.21 rfnmoshv
2059$2059 IOVSS|VSS AVDD|IOVDD \$1143 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2060 r0 *1 4.1,1059.21 rfnmoshv
2060$2060 \$1143 AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2061 r0 *1 4.98,1059.21 rfnmoshv
2061$2061 IOVSS|VSS AVDD|IOVDD \$1143 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2062 r0 *1 5.86,1059.21 rfnmoshv
2062$2062 \$1143 AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2063 r0 *1 6.74,1059.21 rfnmoshv
2063$2063 IOVSS|VSS AVDD|IOVDD \$1143 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2064 r0 *1 7.62,1059.21 rfnmoshv
2064$2064 \$1143 AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2065 r0 *1 13,1059.21 rfnmoshv
2065$2065 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2066 r0 *1 22.88,1059.21 rfnmoshv
2066$2066 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2067 r0 *1 32.76,1059.21 rfnmoshv
2067$2067 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2068 r0 *1 42.64,1059.21 rfnmoshv
2068$2068 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2069 r0 *1 52.52,1059.21 rfnmoshv
2069$2069 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2070 r0 *1 62.4,1059.21 rfnmoshv
2070$2070 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2071 r0 *1 72.28,1059.21 rfnmoshv
2071$2071 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2072 r0 *1 303.22,1059.21 rfnmoshv
2072$2072 IOVSS|VSS IOVDD \$1144 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2073 r0 *1 304.1,1059.21 rfnmoshv
2073$2073 \$1144 IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2074 r0 *1 304.98,1059.21 rfnmoshv
2074$2074 IOVSS|VSS IOVDD \$1144 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2075 r0 *1 305.86,1059.21 rfnmoshv
2075$2075 \$1144 IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2076 r0 *1 306.74,1059.21 rfnmoshv
2076$2076 IOVSS|VSS IOVDD \$1144 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2077 r0 *1 307.62,1059.21 rfnmoshv
2077$2077 \$1144 IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2078 r0 *1 313,1059.21 rfnmoshv
2078$2078 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2079 r0 *1 322.88,1059.21 rfnmoshv
2079$2079 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2080 r0 *1 332.76,1059.21 rfnmoshv
2080$2080 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2081 r0 *1 342.64,1059.21 rfnmoshv
2081$2081 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2082 r0 *1 352.52,1059.21 rfnmoshv
2082$2082 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2083 r0 *1 362.4,1059.21 rfnmoshv
2083$2083 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2084 r0 *1 372.28,1059.21 rfnmoshv
2084$2084 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2085 r0 *1 703.22,1059.21 rfnmoshv
2085$2085 IOVSS|VSS VDD \$1145 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2086 r0 *1 704.1,1059.21 rfnmoshv
2086$2086 \$1145 VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2087 r0 *1 704.98,1059.21 rfnmoshv
2087$2087 IOVSS|VSS VDD \$1145 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2088 r0 *1 705.86,1059.21 rfnmoshv
2088$2088 \$1145 VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2089 r0 *1 706.74,1059.21 rfnmoshv
2089$2089 IOVSS|VSS VDD \$1145 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2090 r0 *1 707.62,1059.21 rfnmoshv
2090$2090 \$1145 VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2091 r0 *1 713,1059.21 rfnmoshv
2091$2091 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2092 r0 *1 722.88,1059.21 rfnmoshv
2092$2092 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2093 r0 *1 732.76,1059.21 rfnmoshv
2093$2093 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2094 r0 *1 742.64,1059.21 rfnmoshv
2094$2094 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2095 r0 *1 752.52,1059.21 rfnmoshv
2095$2095 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2096 r0 *1 762.4,1059.21 rfnmoshv
2096$2096 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2097 r0 *1 772.28,1059.21 rfnmoshv
2097$2097 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2098 r0 *1 3.22,1068.46 rfnmoshv
2098$2098 IOVSS|VSS AVDD|IOVDD \$1143 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2099 r0 *1 4.1,1068.46 rfnmoshv
2099$2099 \$1143 AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2100 r0 *1 4.98,1068.46 rfnmoshv
2100$2100 IOVSS|VSS AVDD|IOVDD \$1143 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2101 r0 *1 5.86,1068.46 rfnmoshv
2101$2101 \$1143 AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2102 r0 *1 6.74,1068.46 rfnmoshv
2102$2102 IOVSS|VSS AVDD|IOVDD \$1143 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2103 r0 *1 7.62,1068.46 rfnmoshv
2103$2103 \$1143 AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2104 r0 *1 13,1068.46 rfnmoshv
2104$2104 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2105 r0 *1 22.88,1068.46 rfnmoshv
2105$2105 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2106 r0 *1 32.76,1068.46 rfnmoshv
2106$2106 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2107 r0 *1 42.64,1068.46 rfnmoshv
2107$2107 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2108 r0 *1 52.52,1068.46 rfnmoshv
2108$2108 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2109 r0 *1 62.4,1068.46 rfnmoshv
2109$2109 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2110 r0 *1 72.28,1068.46 rfnmoshv
2110$2110 IOVSS|VSS AVDD|IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2111 r0 *1 303.22,1068.46 rfnmoshv
2111$2111 IOVSS|VSS IOVDD \$1144 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2112 r0 *1 304.1,1068.46 rfnmoshv
2112$2112 \$1144 IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2113 r0 *1 304.98,1068.46 rfnmoshv
2113$2113 IOVSS|VSS IOVDD \$1144 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2114 r0 *1 305.86,1068.46 rfnmoshv
2114$2114 \$1144 IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2115 r0 *1 306.74,1068.46 rfnmoshv
2115$2115 IOVSS|VSS IOVDD \$1144 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2116 r0 *1 307.62,1068.46 rfnmoshv
2116$2116 \$1144 IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2117 r0 *1 313,1068.46 rfnmoshv
2117$2117 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2118 r0 *1 322.88,1068.46 rfnmoshv
2118$2118 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2119 r0 *1 332.76,1068.46 rfnmoshv
2119$2119 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2120 r0 *1 342.64,1068.46 rfnmoshv
2120$2120 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2121 r0 *1 352.52,1068.46 rfnmoshv
2121$2121 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2122 r0 *1 362.4,1068.46 rfnmoshv
2122$2122 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2123 r0 *1 372.28,1068.46 rfnmoshv
2123$2123 IOVSS|VSS IOVDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2124 r0 *1 703.22,1068.46 rfnmoshv
2124$2124 IOVSS|VSS VDD \$1145 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2125 r0 *1 704.1,1068.46 rfnmoshv
2125$2125 \$1145 VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2126 r0 *1 704.98,1068.46 rfnmoshv
2126$2126 IOVSS|VSS VDD \$1145 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2127 r0 *1 705.86,1068.46 rfnmoshv
2127$2127 \$1145 VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2128 r0 *1 706.74,1068.46 rfnmoshv
2128$2128 IOVSS|VSS VDD \$1145 IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2129 r0 *1 707.62,1068.46 rfnmoshv
2129$2129 \$1145 VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=0.4999999999999999
* device instance $2130 r0 *1 713,1068.46 rfnmoshv
2130$2130 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2131 r0 *1 722.88,1068.46 rfnmoshv
2131$2131 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2132 r0 *1 732.76,1068.46 rfnmoshv
2132$2132 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2133 r0 *1 742.64,1068.46 rfnmoshv
2133$2133 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2134 r0 *1 752.52,1068.46 rfnmoshv
2134$2134 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2135 r0 *1 762.4,1068.46 rfnmoshv
2135$2135 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2136 r0 *1 772.28,1068.46 rfnmoshv
2136$2136 IOVSS|VSS VDD IOVSS|VSS IOVSS|VSS rfnmoshv W=8.999999999999998
+ L=9.499999999999996
* device instance $2137 r0 *1 8.155,1114.53 rfnmoshv
2137$2137 IOVSS|VSS \$1143 \$1316 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2138 r0 *1 9.935,1114.53 rfnmoshv
2138$2138 \$1316 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2139 r0 *1 11.175,1114.53 rfnmoshv
2139$2139 IOVSS|VSS \$1143 \$1317 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2140 r0 *1 12.955,1114.53 rfnmoshv
2140$2140 \$1317 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2141 r0 *1 14.195,1114.53 rfnmoshv
2141$2141 IOVSS|VSS \$1143 \$1318 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2142 r0 *1 15.975,1114.53 rfnmoshv
2142$2142 \$1318 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2143 r0 *1 17.215,1114.53 rfnmoshv
2143$2143 IOVSS|VSS \$1143 \$1319 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2144 r0 *1 18.995,1114.53 rfnmoshv
2144$2144 \$1319 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2145 r0 *1 20.235,1114.53 rfnmoshv
2145$2145 IOVSS|VSS \$1143 \$1320 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2146 r0 *1 22.015,1114.53 rfnmoshv
2146$2146 \$1320 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2147 r0 *1 23.255,1114.53 rfnmoshv
2147$2147 IOVSS|VSS \$1143 \$1321 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2148 r0 *1 25.035,1114.53 rfnmoshv
2148$2148 \$1321 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2149 r0 *1 26.275,1114.53 rfnmoshv
2149$2149 IOVSS|VSS \$1143 \$1322 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2150 r0 *1 28.055,1114.53 rfnmoshv
2150$2150 \$1322 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2151 r0 *1 29.295,1114.53 rfnmoshv
2151$2151 IOVSS|VSS \$1143 \$1323 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2152 r0 *1 31.075,1114.53 rfnmoshv
2152$2152 \$1323 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2153 r0 *1 32.315,1114.53 rfnmoshv
2153$2153 IOVSS|VSS \$1143 \$1324 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2154 r0 *1 34.095,1114.53 rfnmoshv
2154$2154 \$1324 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2155 r0 *1 35.335,1114.53 rfnmoshv
2155$2155 IOVSS|VSS \$1143 \$1325 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2156 r0 *1 37.115,1114.53 rfnmoshv
2156$2156 \$1325 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2157 r0 *1 38.355,1114.53 rfnmoshv
2157$2157 IOVSS|VSS \$1143 \$1326 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2158 r0 *1 40.135,1114.53 rfnmoshv
2158$2158 \$1326 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2159 r0 *1 41.375,1114.53 rfnmoshv
2159$2159 IOVSS|VSS \$1143 \$1327 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2160 r0 *1 43.155,1114.53 rfnmoshv
2160$2160 \$1327 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2161 r0 *1 44.395,1114.53 rfnmoshv
2161$2161 IOVSS|VSS \$1143 \$1328 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2162 r0 *1 46.175,1114.53 rfnmoshv
2162$2162 \$1328 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2163 r0 *1 47.415,1114.53 rfnmoshv
2163$2163 IOVSS|VSS \$1143 \$1329 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2164 r0 *1 49.195,1114.53 rfnmoshv
2164$2164 \$1329 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2165 r0 *1 50.435,1114.53 rfnmoshv
2165$2165 IOVSS|VSS \$1143 \$1330 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2166 r0 *1 52.215,1114.53 rfnmoshv
2166$2166 \$1330 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2167 r0 *1 53.455,1114.53 rfnmoshv
2167$2167 IOVSS|VSS \$1143 \$1331 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2168 r0 *1 55.235,1114.53 rfnmoshv
2168$2168 \$1331 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2169 r0 *1 56.475,1114.53 rfnmoshv
2169$2169 IOVSS|VSS \$1143 \$1332 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2170 r0 *1 58.255,1114.53 rfnmoshv
2170$2170 \$1332 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2171 r0 *1 59.495,1114.53 rfnmoshv
2171$2171 IOVSS|VSS \$1143 \$1333 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2172 r0 *1 61.275,1114.53 rfnmoshv
2172$2172 \$1333 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2173 r0 *1 62.515,1114.53 rfnmoshv
2173$2173 IOVSS|VSS \$1143 \$1334 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2174 r0 *1 64.295,1114.53 rfnmoshv
2174$2174 \$1334 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2175 r0 *1 65.535,1114.53 rfnmoshv
2175$2175 IOVSS|VSS \$1143 \$1335 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2176 r0 *1 67.315,1114.53 rfnmoshv
2176$2176 \$1335 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2177 r0 *1 68.555,1114.53 rfnmoshv
2177$2177 IOVSS|VSS \$1143 \$1336 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2178 r0 *1 70.335,1114.53 rfnmoshv
2178$2178 \$1336 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2179 r0 *1 71.575,1114.53 rfnmoshv
2179$2179 IOVSS|VSS \$1143 \$1337 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2180 r0 *1 308.155,1114.53 rfnmoshv
2180$2180 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2181 r0 *1 309.935,1114.53 rfnmoshv
2181$2181 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2182 r0 *1 311.175,1114.53 rfnmoshv
2182$2182 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2183 r0 *1 312.955,1114.53 rfnmoshv
2183$2183 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2184 r0 *1 314.195,1114.53 rfnmoshv
2184$2184 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2185 r0 *1 315.975,1114.53 rfnmoshv
2185$2185 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2186 r0 *1 317.215,1114.53 rfnmoshv
2186$2186 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2187 r0 *1 318.995,1114.53 rfnmoshv
2187$2187 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2188 r0 *1 320.235,1114.53 rfnmoshv
2188$2188 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2189 r0 *1 322.015,1114.53 rfnmoshv
2189$2189 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2190 r0 *1 323.255,1114.53 rfnmoshv
2190$2190 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2191 r0 *1 325.035,1114.53 rfnmoshv
2191$2191 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2192 r0 *1 326.275,1114.53 rfnmoshv
2192$2192 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2193 r0 *1 328.055,1114.53 rfnmoshv
2193$2193 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2194 r0 *1 329.295,1114.53 rfnmoshv
2194$2194 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2195 r0 *1 331.075,1114.53 rfnmoshv
2195$2195 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2196 r0 *1 332.315,1114.53 rfnmoshv
2196$2196 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2197 r0 *1 334.095,1114.53 rfnmoshv
2197$2197 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2198 r0 *1 335.335,1114.53 rfnmoshv
2198$2198 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2199 r0 *1 337.115,1114.53 rfnmoshv
2199$2199 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2200 r0 *1 338.355,1114.53 rfnmoshv
2200$2200 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2201 r0 *1 340.135,1114.53 rfnmoshv
2201$2201 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2202 r0 *1 341.375,1114.53 rfnmoshv
2202$2202 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2203 r0 *1 343.155,1114.53 rfnmoshv
2203$2203 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2204 r0 *1 344.395,1114.53 rfnmoshv
2204$2204 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2205 r0 *1 346.175,1114.53 rfnmoshv
2205$2205 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2206 r0 *1 347.415,1114.53 rfnmoshv
2206$2206 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2207 r0 *1 349.195,1114.53 rfnmoshv
2207$2207 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2208 r0 *1 350.435,1114.53 rfnmoshv
2208$2208 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2209 r0 *1 352.215,1114.53 rfnmoshv
2209$2209 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2210 r0 *1 353.455,1114.53 rfnmoshv
2210$2210 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2211 r0 *1 355.235,1114.53 rfnmoshv
2211$2211 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2212 r0 *1 356.475,1114.53 rfnmoshv
2212$2212 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2213 r0 *1 358.255,1114.53 rfnmoshv
2213$2213 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2214 r0 *1 359.495,1114.53 rfnmoshv
2214$2214 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2215 r0 *1 361.275,1114.53 rfnmoshv
2215$2215 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2216 r0 *1 362.515,1114.53 rfnmoshv
2216$2216 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2217 r0 *1 364.295,1114.53 rfnmoshv
2217$2217 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2218 r0 *1 365.535,1114.53 rfnmoshv
2218$2218 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2219 r0 *1 367.315,1114.53 rfnmoshv
2219$2219 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2220 r0 *1 368.555,1114.53 rfnmoshv
2220$2220 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2221 r0 *1 370.335,1114.53 rfnmoshv
2221$2221 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2222 r0 *1 371.575,1114.53 rfnmoshv
2222$2222 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2223 r0 *1 708.155,1114.53 rfnmoshv
2223$2223 IOVSS|VSS \$1145 \$1338 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2224 r0 *1 709.935,1114.53 rfnmoshv
2224$2224 \$1338 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2225 r0 *1 711.175,1114.53 rfnmoshv
2225$2225 IOVSS|VSS \$1145 \$1339 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2226 r0 *1 712.955,1114.53 rfnmoshv
2226$2226 \$1339 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2227 r0 *1 714.195,1114.53 rfnmoshv
2227$2227 IOVSS|VSS \$1145 \$1340 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2228 r0 *1 715.975,1114.53 rfnmoshv
2228$2228 \$1340 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2229 r0 *1 717.215,1114.53 rfnmoshv
2229$2229 IOVSS|VSS \$1145 \$1341 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2230 r0 *1 718.995,1114.53 rfnmoshv
2230$2230 \$1341 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2231 r0 *1 720.235,1114.53 rfnmoshv
2231$2231 IOVSS|VSS \$1145 \$1342 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2232 r0 *1 722.015,1114.53 rfnmoshv
2232$2232 \$1342 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2233 r0 *1 723.255,1114.53 rfnmoshv
2233$2233 IOVSS|VSS \$1145 \$1343 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2234 r0 *1 725.035,1114.53 rfnmoshv
2234$2234 \$1343 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2235 r0 *1 726.275,1114.53 rfnmoshv
2235$2235 IOVSS|VSS \$1145 \$1344 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2236 r0 *1 728.055,1114.53 rfnmoshv
2236$2236 \$1344 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2237 r0 *1 729.295,1114.53 rfnmoshv
2237$2237 IOVSS|VSS \$1145 \$1345 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2238 r0 *1 731.075,1114.53 rfnmoshv
2238$2238 \$1345 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2239 r0 *1 732.315,1114.53 rfnmoshv
2239$2239 IOVSS|VSS \$1145 \$1346 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2240 r0 *1 734.095,1114.53 rfnmoshv
2240$2240 \$1346 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2241 r0 *1 735.335,1114.53 rfnmoshv
2241$2241 IOVSS|VSS \$1145 \$1347 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2242 r0 *1 737.115,1114.53 rfnmoshv
2242$2242 \$1347 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2243 r0 *1 738.355,1114.53 rfnmoshv
2243$2243 IOVSS|VSS \$1145 \$1348 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2244 r0 *1 740.135,1114.53 rfnmoshv
2244$2244 \$1348 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2245 r0 *1 741.375,1114.53 rfnmoshv
2245$2245 IOVSS|VSS \$1145 \$1349 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2246 r0 *1 743.155,1114.53 rfnmoshv
2246$2246 \$1349 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2247 r0 *1 744.395,1114.53 rfnmoshv
2247$2247 IOVSS|VSS \$1145 \$1350 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2248 r0 *1 746.175,1114.53 rfnmoshv
2248$2248 \$1350 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2249 r0 *1 747.415,1114.53 rfnmoshv
2249$2249 IOVSS|VSS \$1145 \$1351 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2250 r0 *1 749.195,1114.53 rfnmoshv
2250$2250 \$1351 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2251 r0 *1 750.435,1114.53 rfnmoshv
2251$2251 IOVSS|VSS \$1145 \$1352 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2252 r0 *1 752.215,1114.53 rfnmoshv
2252$2252 \$1352 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2253 r0 *1 753.455,1114.53 rfnmoshv
2253$2253 IOVSS|VSS \$1145 \$1353 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2254 r0 *1 755.235,1114.53 rfnmoshv
2254$2254 \$1353 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2255 r0 *1 756.475,1114.53 rfnmoshv
2255$2255 IOVSS|VSS \$1145 \$1354 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2256 r0 *1 758.255,1114.53 rfnmoshv
2256$2256 \$1354 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2257 r0 *1 759.495,1114.53 rfnmoshv
2257$2257 IOVSS|VSS \$1145 \$1355 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2258 r0 *1 761.275,1114.53 rfnmoshv
2258$2258 \$1355 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2259 r0 *1 762.515,1114.53 rfnmoshv
2259$2259 IOVSS|VSS \$1145 \$1356 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2260 r0 *1 764.295,1114.53 rfnmoshv
2260$2260 \$1356 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2261 r0 *1 765.535,1114.53 rfnmoshv
2261$2261 IOVSS|VSS \$1145 \$1357 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2262 r0 *1 767.315,1114.53 rfnmoshv
2262$2262 \$1357 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2263 r0 *1 768.555,1114.53 rfnmoshv
2263$2263 IOVSS|VSS \$1145 \$1358 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2264 r0 *1 770.335,1114.53 rfnmoshv
2264$2264 \$1358 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2265 r0 *1 771.575,1114.53 rfnmoshv
2265$2265 IOVSS|VSS \$1145 \$1359 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2266 r0 *1 8.155,1119.37 rfnmoshv
2266$2266 IOVSS|VSS \$1143 \$1316 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2267 r0 *1 9.935,1119.37 rfnmoshv
2267$2267 \$1316 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2268 r0 *1 11.175,1119.37 rfnmoshv
2268$2268 IOVSS|VSS \$1143 \$1317 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2269 r0 *1 12.955,1119.37 rfnmoshv
2269$2269 \$1317 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2270 r0 *1 14.195,1119.37 rfnmoshv
2270$2270 IOVSS|VSS \$1143 \$1318 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2271 r0 *1 15.975,1119.37 rfnmoshv
2271$2271 \$1318 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2272 r0 *1 17.215,1119.37 rfnmoshv
2272$2272 IOVSS|VSS \$1143 \$1319 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2273 r0 *1 18.995,1119.37 rfnmoshv
2273$2273 \$1319 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2274 r0 *1 20.235,1119.37 rfnmoshv
2274$2274 IOVSS|VSS \$1143 \$1320 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2275 r0 *1 22.015,1119.37 rfnmoshv
2275$2275 \$1320 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2276 r0 *1 23.255,1119.37 rfnmoshv
2276$2276 IOVSS|VSS \$1143 \$1321 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2277 r0 *1 25.035,1119.37 rfnmoshv
2277$2277 \$1321 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2278 r0 *1 26.275,1119.37 rfnmoshv
2278$2278 IOVSS|VSS \$1143 \$1322 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2279 r0 *1 28.055,1119.37 rfnmoshv
2279$2279 \$1322 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2280 r0 *1 29.295,1119.37 rfnmoshv
2280$2280 IOVSS|VSS \$1143 \$1323 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2281 r0 *1 31.075,1119.37 rfnmoshv
2281$2281 \$1323 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2282 r0 *1 32.315,1119.37 rfnmoshv
2282$2282 IOVSS|VSS \$1143 \$1324 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2283 r0 *1 34.095,1119.37 rfnmoshv
2283$2283 \$1324 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2284 r0 *1 35.335,1119.37 rfnmoshv
2284$2284 IOVSS|VSS \$1143 \$1325 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2285 r0 *1 37.115,1119.37 rfnmoshv
2285$2285 \$1325 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2286 r0 *1 38.355,1119.37 rfnmoshv
2286$2286 IOVSS|VSS \$1143 \$1326 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2287 r0 *1 40.135,1119.37 rfnmoshv
2287$2287 \$1326 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2288 r0 *1 41.375,1119.37 rfnmoshv
2288$2288 IOVSS|VSS \$1143 \$1327 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2289 r0 *1 43.155,1119.37 rfnmoshv
2289$2289 \$1327 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2290 r0 *1 44.395,1119.37 rfnmoshv
2290$2290 IOVSS|VSS \$1143 \$1328 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2291 r0 *1 46.175,1119.37 rfnmoshv
2291$2291 \$1328 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2292 r0 *1 47.415,1119.37 rfnmoshv
2292$2292 IOVSS|VSS \$1143 \$1329 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2293 r0 *1 49.195,1119.37 rfnmoshv
2293$2293 \$1329 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2294 r0 *1 50.435,1119.37 rfnmoshv
2294$2294 IOVSS|VSS \$1143 \$1330 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2295 r0 *1 52.215,1119.37 rfnmoshv
2295$2295 \$1330 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2296 r0 *1 53.455,1119.37 rfnmoshv
2296$2296 IOVSS|VSS \$1143 \$1331 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2297 r0 *1 55.235,1119.37 rfnmoshv
2297$2297 \$1331 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2298 r0 *1 56.475,1119.37 rfnmoshv
2298$2298 IOVSS|VSS \$1143 \$1332 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2299 r0 *1 58.255,1119.37 rfnmoshv
2299$2299 \$1332 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2300 r0 *1 59.495,1119.37 rfnmoshv
2300$2300 IOVSS|VSS \$1143 \$1333 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2301 r0 *1 61.275,1119.37 rfnmoshv
2301$2301 \$1333 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2302 r0 *1 62.515,1119.37 rfnmoshv
2302$2302 IOVSS|VSS \$1143 \$1334 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2303 r0 *1 64.295,1119.37 rfnmoshv
2303$2303 \$1334 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2304 r0 *1 65.535,1119.37 rfnmoshv
2304$2304 IOVSS|VSS \$1143 \$1335 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2305 r0 *1 67.315,1119.37 rfnmoshv
2305$2305 \$1335 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2306 r0 *1 68.555,1119.37 rfnmoshv
2306$2306 IOVSS|VSS \$1143 \$1336 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2307 r0 *1 70.335,1119.37 rfnmoshv
2307$2307 \$1336 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2308 r0 *1 71.575,1119.37 rfnmoshv
2308$2308 IOVSS|VSS \$1143 \$1337 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2309 r0 *1 308.155,1119.37 rfnmoshv
2309$2309 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2310 r0 *1 309.935,1119.37 rfnmoshv
2310$2310 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2311 r0 *1 311.175,1119.37 rfnmoshv
2311$2311 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2312 r0 *1 312.955,1119.37 rfnmoshv
2312$2312 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2313 r0 *1 314.195,1119.37 rfnmoshv
2313$2313 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2314 r0 *1 315.975,1119.37 rfnmoshv
2314$2314 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2315 r0 *1 317.215,1119.37 rfnmoshv
2315$2315 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2316 r0 *1 318.995,1119.37 rfnmoshv
2316$2316 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2317 r0 *1 320.235,1119.37 rfnmoshv
2317$2317 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2318 r0 *1 322.015,1119.37 rfnmoshv
2318$2318 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2319 r0 *1 323.255,1119.37 rfnmoshv
2319$2319 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2320 r0 *1 325.035,1119.37 rfnmoshv
2320$2320 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2321 r0 *1 326.275,1119.37 rfnmoshv
2321$2321 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2322 r0 *1 328.055,1119.37 rfnmoshv
2322$2322 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2323 r0 *1 329.295,1119.37 rfnmoshv
2323$2323 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2324 r0 *1 331.075,1119.37 rfnmoshv
2324$2324 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2325 r0 *1 332.315,1119.37 rfnmoshv
2325$2325 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2326 r0 *1 334.095,1119.37 rfnmoshv
2326$2326 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2327 r0 *1 335.335,1119.37 rfnmoshv
2327$2327 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2328 r0 *1 337.115,1119.37 rfnmoshv
2328$2328 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2329 r0 *1 338.355,1119.37 rfnmoshv
2329$2329 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2330 r0 *1 340.135,1119.37 rfnmoshv
2330$2330 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2331 r0 *1 341.375,1119.37 rfnmoshv
2331$2331 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2332 r0 *1 343.155,1119.37 rfnmoshv
2332$2332 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2333 r0 *1 344.395,1119.37 rfnmoshv
2333$2333 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2334 r0 *1 346.175,1119.37 rfnmoshv
2334$2334 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2335 r0 *1 347.415,1119.37 rfnmoshv
2335$2335 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2336 r0 *1 349.195,1119.37 rfnmoshv
2336$2336 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2337 r0 *1 350.435,1119.37 rfnmoshv
2337$2337 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2338 r0 *1 352.215,1119.37 rfnmoshv
2338$2338 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2339 r0 *1 353.455,1119.37 rfnmoshv
2339$2339 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2340 r0 *1 355.235,1119.37 rfnmoshv
2340$2340 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2341 r0 *1 356.475,1119.37 rfnmoshv
2341$2341 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2342 r0 *1 358.255,1119.37 rfnmoshv
2342$2342 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2343 r0 *1 359.495,1119.37 rfnmoshv
2343$2343 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2344 r0 *1 361.275,1119.37 rfnmoshv
2344$2344 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2345 r0 *1 362.515,1119.37 rfnmoshv
2345$2345 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2346 r0 *1 364.295,1119.37 rfnmoshv
2346$2346 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2347 r0 *1 365.535,1119.37 rfnmoshv
2347$2347 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2348 r0 *1 367.315,1119.37 rfnmoshv
2348$2348 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2349 r0 *1 368.555,1119.37 rfnmoshv
2349$2349 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2350 r0 *1 370.335,1119.37 rfnmoshv
2350$2350 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2351 r0 *1 371.575,1119.37 rfnmoshv
2351$2351 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2352 r0 *1 708.155,1119.37 rfnmoshv
2352$2352 IOVSS|VSS \$1145 \$1338 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2353 r0 *1 709.935,1119.37 rfnmoshv
2353$2353 \$1338 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2354 r0 *1 711.175,1119.37 rfnmoshv
2354$2354 IOVSS|VSS \$1145 \$1339 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2355 r0 *1 712.955,1119.37 rfnmoshv
2355$2355 \$1339 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2356 r0 *1 714.195,1119.37 rfnmoshv
2356$2356 IOVSS|VSS \$1145 \$1340 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2357 r0 *1 715.975,1119.37 rfnmoshv
2357$2357 \$1340 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2358 r0 *1 717.215,1119.37 rfnmoshv
2358$2358 IOVSS|VSS \$1145 \$1341 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2359 r0 *1 718.995,1119.37 rfnmoshv
2359$2359 \$1341 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2360 r0 *1 720.235,1119.37 rfnmoshv
2360$2360 IOVSS|VSS \$1145 \$1342 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2361 r0 *1 722.015,1119.37 rfnmoshv
2361$2361 \$1342 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2362 r0 *1 723.255,1119.37 rfnmoshv
2362$2362 IOVSS|VSS \$1145 \$1343 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2363 r0 *1 725.035,1119.37 rfnmoshv
2363$2363 \$1343 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2364 r0 *1 726.275,1119.37 rfnmoshv
2364$2364 IOVSS|VSS \$1145 \$1344 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2365 r0 *1 728.055,1119.37 rfnmoshv
2365$2365 \$1344 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2366 r0 *1 729.295,1119.37 rfnmoshv
2366$2366 IOVSS|VSS \$1145 \$1345 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2367 r0 *1 731.075,1119.37 rfnmoshv
2367$2367 \$1345 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2368 r0 *1 732.315,1119.37 rfnmoshv
2368$2368 IOVSS|VSS \$1145 \$1346 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2369 r0 *1 734.095,1119.37 rfnmoshv
2369$2369 \$1346 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2370 r0 *1 735.335,1119.37 rfnmoshv
2370$2370 IOVSS|VSS \$1145 \$1347 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2371 r0 *1 737.115,1119.37 rfnmoshv
2371$2371 \$1347 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2372 r0 *1 738.355,1119.37 rfnmoshv
2372$2372 IOVSS|VSS \$1145 \$1348 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2373 r0 *1 740.135,1119.37 rfnmoshv
2373$2373 \$1348 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2374 r0 *1 741.375,1119.37 rfnmoshv
2374$2374 IOVSS|VSS \$1145 \$1349 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2375 r0 *1 743.155,1119.37 rfnmoshv
2375$2375 \$1349 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2376 r0 *1 744.395,1119.37 rfnmoshv
2376$2376 IOVSS|VSS \$1145 \$1350 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2377 r0 *1 746.175,1119.37 rfnmoshv
2377$2377 \$1350 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2378 r0 *1 747.415,1119.37 rfnmoshv
2378$2378 IOVSS|VSS \$1145 \$1351 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2379 r0 *1 749.195,1119.37 rfnmoshv
2379$2379 \$1351 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2380 r0 *1 750.435,1119.37 rfnmoshv
2380$2380 IOVSS|VSS \$1145 \$1352 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2381 r0 *1 752.215,1119.37 rfnmoshv
2381$2381 \$1352 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2382 r0 *1 753.455,1119.37 rfnmoshv
2382$2382 IOVSS|VSS \$1145 \$1353 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2383 r0 *1 755.235,1119.37 rfnmoshv
2383$2383 \$1353 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2384 r0 *1 756.475,1119.37 rfnmoshv
2384$2384 IOVSS|VSS \$1145 \$1354 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2385 r0 *1 758.255,1119.37 rfnmoshv
2385$2385 \$1354 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2386 r0 *1 759.495,1119.37 rfnmoshv
2386$2386 IOVSS|VSS \$1145 \$1355 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2387 r0 *1 761.275,1119.37 rfnmoshv
2387$2387 \$1355 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2388 r0 *1 762.515,1119.37 rfnmoshv
2388$2388 IOVSS|VSS \$1145 \$1356 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2389 r0 *1 764.295,1119.37 rfnmoshv
2389$2389 \$1356 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2390 r0 *1 765.535,1119.37 rfnmoshv
2390$2390 IOVSS|VSS \$1145 \$1357 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2391 r0 *1 767.315,1119.37 rfnmoshv
2391$2391 \$1357 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2392 r0 *1 768.555,1119.37 rfnmoshv
2392$2392 IOVSS|VSS \$1145 \$1358 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2393 r0 *1 770.335,1119.37 rfnmoshv
2393$2393 \$1358 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2394 r0 *1 771.575,1119.37 rfnmoshv
2394$2394 IOVSS|VSS \$1145 \$1359 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2395 r0 *1 8.155,1124.21 rfnmoshv
2395$2395 IOVSS|VSS \$1143 \$1316 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2396 r0 *1 9.935,1124.21 rfnmoshv
2396$2396 \$1316 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2397 r0 *1 11.175,1124.21 rfnmoshv
2397$2397 IOVSS|VSS \$1143 \$1317 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2398 r0 *1 12.955,1124.21 rfnmoshv
2398$2398 \$1317 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2399 r0 *1 14.195,1124.21 rfnmoshv
2399$2399 IOVSS|VSS \$1143 \$1318 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2400 r0 *1 15.975,1124.21 rfnmoshv
2400$2400 \$1318 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2401 r0 *1 17.215,1124.21 rfnmoshv
2401$2401 IOVSS|VSS \$1143 \$1319 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2402 r0 *1 18.995,1124.21 rfnmoshv
2402$2402 \$1319 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2403 r0 *1 20.235,1124.21 rfnmoshv
2403$2403 IOVSS|VSS \$1143 \$1320 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2404 r0 *1 22.015,1124.21 rfnmoshv
2404$2404 \$1320 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2405 r0 *1 23.255,1124.21 rfnmoshv
2405$2405 IOVSS|VSS \$1143 \$1321 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2406 r0 *1 25.035,1124.21 rfnmoshv
2406$2406 \$1321 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2407 r0 *1 26.275,1124.21 rfnmoshv
2407$2407 IOVSS|VSS \$1143 \$1322 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2408 r0 *1 28.055,1124.21 rfnmoshv
2408$2408 \$1322 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2409 r0 *1 29.295,1124.21 rfnmoshv
2409$2409 IOVSS|VSS \$1143 \$1323 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2410 r0 *1 31.075,1124.21 rfnmoshv
2410$2410 \$1323 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2411 r0 *1 32.315,1124.21 rfnmoshv
2411$2411 IOVSS|VSS \$1143 \$1324 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2412 r0 *1 34.095,1124.21 rfnmoshv
2412$2412 \$1324 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2413 r0 *1 35.335,1124.21 rfnmoshv
2413$2413 IOVSS|VSS \$1143 \$1325 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2414 r0 *1 37.115,1124.21 rfnmoshv
2414$2414 \$1325 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2415 r0 *1 38.355,1124.21 rfnmoshv
2415$2415 IOVSS|VSS \$1143 \$1326 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2416 r0 *1 40.135,1124.21 rfnmoshv
2416$2416 \$1326 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2417 r0 *1 41.375,1124.21 rfnmoshv
2417$2417 IOVSS|VSS \$1143 \$1327 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2418 r0 *1 43.155,1124.21 rfnmoshv
2418$2418 \$1327 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2419 r0 *1 44.395,1124.21 rfnmoshv
2419$2419 IOVSS|VSS \$1143 \$1328 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2420 r0 *1 46.175,1124.21 rfnmoshv
2420$2420 \$1328 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2421 r0 *1 47.415,1124.21 rfnmoshv
2421$2421 IOVSS|VSS \$1143 \$1329 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2422 r0 *1 49.195,1124.21 rfnmoshv
2422$2422 \$1329 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2423 r0 *1 50.435,1124.21 rfnmoshv
2423$2423 IOVSS|VSS \$1143 \$1330 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2424 r0 *1 52.215,1124.21 rfnmoshv
2424$2424 \$1330 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2425 r0 *1 53.455,1124.21 rfnmoshv
2425$2425 IOVSS|VSS \$1143 \$1331 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2426 r0 *1 55.235,1124.21 rfnmoshv
2426$2426 \$1331 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2427 r0 *1 56.475,1124.21 rfnmoshv
2427$2427 IOVSS|VSS \$1143 \$1332 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2428 r0 *1 58.255,1124.21 rfnmoshv
2428$2428 \$1332 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2429 r0 *1 59.495,1124.21 rfnmoshv
2429$2429 IOVSS|VSS \$1143 \$1333 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2430 r0 *1 61.275,1124.21 rfnmoshv
2430$2430 \$1333 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2431 r0 *1 62.515,1124.21 rfnmoshv
2431$2431 IOVSS|VSS \$1143 \$1334 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2432 r0 *1 64.295,1124.21 rfnmoshv
2432$2432 \$1334 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2433 r0 *1 65.535,1124.21 rfnmoshv
2433$2433 IOVSS|VSS \$1143 \$1335 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2434 r0 *1 67.315,1124.21 rfnmoshv
2434$2434 \$1335 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2435 r0 *1 68.555,1124.21 rfnmoshv
2435$2435 IOVSS|VSS \$1143 \$1336 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2436 r0 *1 70.335,1124.21 rfnmoshv
2436$2436 \$1336 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2437 r0 *1 71.575,1124.21 rfnmoshv
2437$2437 IOVSS|VSS \$1143 \$1337 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2438 r0 *1 308.155,1124.21 rfnmoshv
2438$2438 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2439 r0 *1 309.935,1124.21 rfnmoshv
2439$2439 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2440 r0 *1 311.175,1124.21 rfnmoshv
2440$2440 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2441 r0 *1 312.955,1124.21 rfnmoshv
2441$2441 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2442 r0 *1 314.195,1124.21 rfnmoshv
2442$2442 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2443 r0 *1 315.975,1124.21 rfnmoshv
2443$2443 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2444 r0 *1 317.215,1124.21 rfnmoshv
2444$2444 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2445 r0 *1 318.995,1124.21 rfnmoshv
2445$2445 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2446 r0 *1 320.235,1124.21 rfnmoshv
2446$2446 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2447 r0 *1 322.015,1124.21 rfnmoshv
2447$2447 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2448 r0 *1 323.255,1124.21 rfnmoshv
2448$2448 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2449 r0 *1 325.035,1124.21 rfnmoshv
2449$2449 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2450 r0 *1 326.275,1124.21 rfnmoshv
2450$2450 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2451 r0 *1 328.055,1124.21 rfnmoshv
2451$2451 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2452 r0 *1 329.295,1124.21 rfnmoshv
2452$2452 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2453 r0 *1 331.075,1124.21 rfnmoshv
2453$2453 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2454 r0 *1 332.315,1124.21 rfnmoshv
2454$2454 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2455 r0 *1 334.095,1124.21 rfnmoshv
2455$2455 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2456 r0 *1 335.335,1124.21 rfnmoshv
2456$2456 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2457 r0 *1 337.115,1124.21 rfnmoshv
2457$2457 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2458 r0 *1 338.355,1124.21 rfnmoshv
2458$2458 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2459 r0 *1 340.135,1124.21 rfnmoshv
2459$2459 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2460 r0 *1 341.375,1124.21 rfnmoshv
2460$2460 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2461 r0 *1 343.155,1124.21 rfnmoshv
2461$2461 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2462 r0 *1 344.395,1124.21 rfnmoshv
2462$2462 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2463 r0 *1 346.175,1124.21 rfnmoshv
2463$2463 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2464 r0 *1 347.415,1124.21 rfnmoshv
2464$2464 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2465 r0 *1 349.195,1124.21 rfnmoshv
2465$2465 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2466 r0 *1 350.435,1124.21 rfnmoshv
2466$2466 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2467 r0 *1 352.215,1124.21 rfnmoshv
2467$2467 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2468 r0 *1 353.455,1124.21 rfnmoshv
2468$2468 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2469 r0 *1 355.235,1124.21 rfnmoshv
2469$2469 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2470 r0 *1 356.475,1124.21 rfnmoshv
2470$2470 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2471 r0 *1 358.255,1124.21 rfnmoshv
2471$2471 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2472 r0 *1 359.495,1124.21 rfnmoshv
2472$2472 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2473 r0 *1 361.275,1124.21 rfnmoshv
2473$2473 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2474 r0 *1 362.515,1124.21 rfnmoshv
2474$2474 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2475 r0 *1 364.295,1124.21 rfnmoshv
2475$2475 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2476 r0 *1 365.535,1124.21 rfnmoshv
2476$2476 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2477 r0 *1 367.315,1124.21 rfnmoshv
2477$2477 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2478 r0 *1 368.555,1124.21 rfnmoshv
2478$2478 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2479 r0 *1 370.335,1124.21 rfnmoshv
2479$2479 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2480 r0 *1 371.575,1124.21 rfnmoshv
2480$2480 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2481 r0 *1 708.155,1124.21 rfnmoshv
2481$2481 IOVSS|VSS \$1145 \$1338 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2482 r0 *1 709.935,1124.21 rfnmoshv
2482$2482 \$1338 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2483 r0 *1 711.175,1124.21 rfnmoshv
2483$2483 IOVSS|VSS \$1145 \$1339 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2484 r0 *1 712.955,1124.21 rfnmoshv
2484$2484 \$1339 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2485 r0 *1 714.195,1124.21 rfnmoshv
2485$2485 IOVSS|VSS \$1145 \$1340 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2486 r0 *1 715.975,1124.21 rfnmoshv
2486$2486 \$1340 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2487 r0 *1 717.215,1124.21 rfnmoshv
2487$2487 IOVSS|VSS \$1145 \$1341 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2488 r0 *1 718.995,1124.21 rfnmoshv
2488$2488 \$1341 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2489 r0 *1 720.235,1124.21 rfnmoshv
2489$2489 IOVSS|VSS \$1145 \$1342 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2490 r0 *1 722.015,1124.21 rfnmoshv
2490$2490 \$1342 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2491 r0 *1 723.255,1124.21 rfnmoshv
2491$2491 IOVSS|VSS \$1145 \$1343 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2492 r0 *1 725.035,1124.21 rfnmoshv
2492$2492 \$1343 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2493 r0 *1 726.275,1124.21 rfnmoshv
2493$2493 IOVSS|VSS \$1145 \$1344 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2494 r0 *1 728.055,1124.21 rfnmoshv
2494$2494 \$1344 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2495 r0 *1 729.295,1124.21 rfnmoshv
2495$2495 IOVSS|VSS \$1145 \$1345 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2496 r0 *1 731.075,1124.21 rfnmoshv
2496$2496 \$1345 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2497 r0 *1 732.315,1124.21 rfnmoshv
2497$2497 IOVSS|VSS \$1145 \$1346 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2498 r0 *1 734.095,1124.21 rfnmoshv
2498$2498 \$1346 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2499 r0 *1 735.335,1124.21 rfnmoshv
2499$2499 IOVSS|VSS \$1145 \$1347 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2500 r0 *1 737.115,1124.21 rfnmoshv
2500$2500 \$1347 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2501 r0 *1 738.355,1124.21 rfnmoshv
2501$2501 IOVSS|VSS \$1145 \$1348 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2502 r0 *1 740.135,1124.21 rfnmoshv
2502$2502 \$1348 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2503 r0 *1 741.375,1124.21 rfnmoshv
2503$2503 IOVSS|VSS \$1145 \$1349 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2504 r0 *1 743.155,1124.21 rfnmoshv
2504$2504 \$1349 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2505 r0 *1 744.395,1124.21 rfnmoshv
2505$2505 IOVSS|VSS \$1145 \$1350 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2506 r0 *1 746.175,1124.21 rfnmoshv
2506$2506 \$1350 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2507 r0 *1 747.415,1124.21 rfnmoshv
2507$2507 IOVSS|VSS \$1145 \$1351 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2508 r0 *1 749.195,1124.21 rfnmoshv
2508$2508 \$1351 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2509 r0 *1 750.435,1124.21 rfnmoshv
2509$2509 IOVSS|VSS \$1145 \$1352 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2510 r0 *1 752.215,1124.21 rfnmoshv
2510$2510 \$1352 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2511 r0 *1 753.455,1124.21 rfnmoshv
2511$2511 IOVSS|VSS \$1145 \$1353 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2512 r0 *1 755.235,1124.21 rfnmoshv
2512$2512 \$1353 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2513 r0 *1 756.475,1124.21 rfnmoshv
2513$2513 IOVSS|VSS \$1145 \$1354 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2514 r0 *1 758.255,1124.21 rfnmoshv
2514$2514 \$1354 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2515 r0 *1 759.495,1124.21 rfnmoshv
2515$2515 IOVSS|VSS \$1145 \$1355 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2516 r0 *1 761.275,1124.21 rfnmoshv
2516$2516 \$1355 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2517 r0 *1 762.515,1124.21 rfnmoshv
2517$2517 IOVSS|VSS \$1145 \$1356 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2518 r0 *1 764.295,1124.21 rfnmoshv
2518$2518 \$1356 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2519 r0 *1 765.535,1124.21 rfnmoshv
2519$2519 IOVSS|VSS \$1145 \$1357 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2520 r0 *1 767.315,1124.21 rfnmoshv
2520$2520 \$1357 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2521 r0 *1 768.555,1124.21 rfnmoshv
2521$2521 IOVSS|VSS \$1145 \$1358 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2522 r0 *1 770.335,1124.21 rfnmoshv
2522$2522 \$1358 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2523 r0 *1 771.575,1124.21 rfnmoshv
2523$2523 IOVSS|VSS \$1145 \$1359 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2524 r0 *1 8.155,1129.05 rfnmoshv
2524$2524 IOVSS|VSS \$1143 \$1316 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2525 r0 *1 9.935,1129.05 rfnmoshv
2525$2525 \$1316 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2526 r0 *1 11.175,1129.05 rfnmoshv
2526$2526 IOVSS|VSS \$1143 \$1317 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2527 r0 *1 12.955,1129.05 rfnmoshv
2527$2527 \$1317 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2528 r0 *1 14.195,1129.05 rfnmoshv
2528$2528 IOVSS|VSS \$1143 \$1318 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2529 r0 *1 15.975,1129.05 rfnmoshv
2529$2529 \$1318 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2530 r0 *1 17.215,1129.05 rfnmoshv
2530$2530 IOVSS|VSS \$1143 \$1319 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2531 r0 *1 18.995,1129.05 rfnmoshv
2531$2531 \$1319 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2532 r0 *1 20.235,1129.05 rfnmoshv
2532$2532 IOVSS|VSS \$1143 \$1320 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2533 r0 *1 22.015,1129.05 rfnmoshv
2533$2533 \$1320 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2534 r0 *1 23.255,1129.05 rfnmoshv
2534$2534 IOVSS|VSS \$1143 \$1321 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2535 r0 *1 25.035,1129.05 rfnmoshv
2535$2535 \$1321 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2536 r0 *1 26.275,1129.05 rfnmoshv
2536$2536 IOVSS|VSS \$1143 \$1322 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2537 r0 *1 28.055,1129.05 rfnmoshv
2537$2537 \$1322 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2538 r0 *1 29.295,1129.05 rfnmoshv
2538$2538 IOVSS|VSS \$1143 \$1323 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2539 r0 *1 31.075,1129.05 rfnmoshv
2539$2539 \$1323 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2540 r0 *1 32.315,1129.05 rfnmoshv
2540$2540 IOVSS|VSS \$1143 \$1324 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2541 r0 *1 34.095,1129.05 rfnmoshv
2541$2541 \$1324 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2542 r0 *1 35.335,1129.05 rfnmoshv
2542$2542 IOVSS|VSS \$1143 \$1325 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2543 r0 *1 37.115,1129.05 rfnmoshv
2543$2543 \$1325 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2544 r0 *1 38.355,1129.05 rfnmoshv
2544$2544 IOVSS|VSS \$1143 \$1326 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2545 r0 *1 40.135,1129.05 rfnmoshv
2545$2545 \$1326 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2546 r0 *1 41.375,1129.05 rfnmoshv
2546$2546 IOVSS|VSS \$1143 \$1327 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2547 r0 *1 43.155,1129.05 rfnmoshv
2547$2547 \$1327 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2548 r0 *1 44.395,1129.05 rfnmoshv
2548$2548 IOVSS|VSS \$1143 \$1328 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2549 r0 *1 46.175,1129.05 rfnmoshv
2549$2549 \$1328 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2550 r0 *1 47.415,1129.05 rfnmoshv
2550$2550 IOVSS|VSS \$1143 \$1329 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2551 r0 *1 49.195,1129.05 rfnmoshv
2551$2551 \$1329 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2552 r0 *1 50.435,1129.05 rfnmoshv
2552$2552 IOVSS|VSS \$1143 \$1330 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2553 r0 *1 52.215,1129.05 rfnmoshv
2553$2553 \$1330 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2554 r0 *1 53.455,1129.05 rfnmoshv
2554$2554 IOVSS|VSS \$1143 \$1331 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2555 r0 *1 55.235,1129.05 rfnmoshv
2555$2555 \$1331 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2556 r0 *1 56.475,1129.05 rfnmoshv
2556$2556 IOVSS|VSS \$1143 \$1332 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2557 r0 *1 58.255,1129.05 rfnmoshv
2557$2557 \$1332 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2558 r0 *1 59.495,1129.05 rfnmoshv
2558$2558 IOVSS|VSS \$1143 \$1333 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2559 r0 *1 61.275,1129.05 rfnmoshv
2559$2559 \$1333 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2560 r0 *1 62.515,1129.05 rfnmoshv
2560$2560 IOVSS|VSS \$1143 \$1334 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2561 r0 *1 64.295,1129.05 rfnmoshv
2561$2561 \$1334 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2562 r0 *1 65.535,1129.05 rfnmoshv
2562$2562 IOVSS|VSS \$1143 \$1335 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2563 r0 *1 67.315,1129.05 rfnmoshv
2563$2563 \$1335 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2564 r0 *1 68.555,1129.05 rfnmoshv
2564$2564 IOVSS|VSS \$1143 \$1336 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2565 r0 *1 70.335,1129.05 rfnmoshv
2565$2565 \$1336 \$1143 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2566 r0 *1 71.575,1129.05 rfnmoshv
2566$2566 IOVSS|VSS \$1143 \$1337 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2567 r0 *1 308.155,1129.05 rfnmoshv
2567$2567 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2568 r0 *1 309.935,1129.05 rfnmoshv
2568$2568 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2569 r0 *1 311.175,1129.05 rfnmoshv
2569$2569 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2570 r0 *1 312.955,1129.05 rfnmoshv
2570$2570 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2571 r0 *1 314.195,1129.05 rfnmoshv
2571$2571 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2572 r0 *1 315.975,1129.05 rfnmoshv
2572$2572 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2573 r0 *1 317.215,1129.05 rfnmoshv
2573$2573 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2574 r0 *1 318.995,1129.05 rfnmoshv
2574$2574 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2575 r0 *1 320.235,1129.05 rfnmoshv
2575$2575 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2576 r0 *1 322.015,1129.05 rfnmoshv
2576$2576 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2577 r0 *1 323.255,1129.05 rfnmoshv
2577$2577 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2578 r0 *1 325.035,1129.05 rfnmoshv
2578$2578 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2579 r0 *1 326.275,1129.05 rfnmoshv
2579$2579 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2580 r0 *1 328.055,1129.05 rfnmoshv
2580$2580 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2581 r0 *1 329.295,1129.05 rfnmoshv
2581$2581 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2582 r0 *1 331.075,1129.05 rfnmoshv
2582$2582 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2583 r0 *1 332.315,1129.05 rfnmoshv
2583$2583 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2584 r0 *1 334.095,1129.05 rfnmoshv
2584$2584 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2585 r0 *1 335.335,1129.05 rfnmoshv
2585$2585 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2586 r0 *1 337.115,1129.05 rfnmoshv
2586$2586 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2587 r0 *1 338.355,1129.05 rfnmoshv
2587$2587 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2588 r0 *1 340.135,1129.05 rfnmoshv
2588$2588 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2589 r0 *1 341.375,1129.05 rfnmoshv
2589$2589 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2590 r0 *1 343.155,1129.05 rfnmoshv
2590$2590 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2591 r0 *1 344.395,1129.05 rfnmoshv
2591$2591 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2592 r0 *1 346.175,1129.05 rfnmoshv
2592$2592 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2593 r0 *1 347.415,1129.05 rfnmoshv
2593$2593 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2594 r0 *1 349.195,1129.05 rfnmoshv
2594$2594 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2595 r0 *1 350.435,1129.05 rfnmoshv
2595$2595 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2596 r0 *1 352.215,1129.05 rfnmoshv
2596$2596 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2597 r0 *1 353.455,1129.05 rfnmoshv
2597$2597 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2598 r0 *1 355.235,1129.05 rfnmoshv
2598$2598 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2599 r0 *1 356.475,1129.05 rfnmoshv
2599$2599 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2600 r0 *1 358.255,1129.05 rfnmoshv
2600$2600 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2601 r0 *1 359.495,1129.05 rfnmoshv
2601$2601 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2602 r0 *1 361.275,1129.05 rfnmoshv
2602$2602 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2603 r0 *1 362.515,1129.05 rfnmoshv
2603$2603 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2604 r0 *1 364.295,1129.05 rfnmoshv
2604$2604 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2605 r0 *1 365.535,1129.05 rfnmoshv
2605$2605 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2606 r0 *1 367.315,1129.05 rfnmoshv
2606$2606 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2607 r0 *1 368.555,1129.05 rfnmoshv
2607$2607 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2608 r0 *1 370.335,1129.05 rfnmoshv
2608$2608 IOVDD \$1144 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2609 r0 *1 371.575,1129.05 rfnmoshv
2609$2609 IOVSS|VSS \$1144 IOVDD IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2610 r0 *1 708.155,1129.05 rfnmoshv
2610$2610 IOVSS|VSS \$1145 \$1338 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2611 r0 *1 709.935,1129.05 rfnmoshv
2611$2611 \$1338 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2612 r0 *1 711.175,1129.05 rfnmoshv
2612$2612 IOVSS|VSS \$1145 \$1339 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2613 r0 *1 712.955,1129.05 rfnmoshv
2613$2613 \$1339 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2614 r0 *1 714.195,1129.05 rfnmoshv
2614$2614 IOVSS|VSS \$1145 \$1340 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2615 r0 *1 715.975,1129.05 rfnmoshv
2615$2615 \$1340 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2616 r0 *1 717.215,1129.05 rfnmoshv
2616$2616 IOVSS|VSS \$1145 \$1341 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2617 r0 *1 718.995,1129.05 rfnmoshv
2617$2617 \$1341 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2618 r0 *1 720.235,1129.05 rfnmoshv
2618$2618 IOVSS|VSS \$1145 \$1342 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2619 r0 *1 722.015,1129.05 rfnmoshv
2619$2619 \$1342 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2620 r0 *1 723.255,1129.05 rfnmoshv
2620$2620 IOVSS|VSS \$1145 \$1343 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2621 r0 *1 725.035,1129.05 rfnmoshv
2621$2621 \$1343 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2622 r0 *1 726.275,1129.05 rfnmoshv
2622$2622 IOVSS|VSS \$1145 \$1344 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2623 r0 *1 728.055,1129.05 rfnmoshv
2623$2623 \$1344 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2624 r0 *1 729.295,1129.05 rfnmoshv
2624$2624 IOVSS|VSS \$1145 \$1345 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2625 r0 *1 731.075,1129.05 rfnmoshv
2625$2625 \$1345 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2626 r0 *1 732.315,1129.05 rfnmoshv
2626$2626 IOVSS|VSS \$1145 \$1346 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2627 r0 *1 734.095,1129.05 rfnmoshv
2627$2627 \$1346 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2628 r0 *1 735.335,1129.05 rfnmoshv
2628$2628 IOVSS|VSS \$1145 \$1347 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2629 r0 *1 737.115,1129.05 rfnmoshv
2629$2629 \$1347 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2630 r0 *1 738.355,1129.05 rfnmoshv
2630$2630 IOVSS|VSS \$1145 \$1348 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2631 r0 *1 740.135,1129.05 rfnmoshv
2631$2631 \$1348 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2632 r0 *1 741.375,1129.05 rfnmoshv
2632$2632 IOVSS|VSS \$1145 \$1349 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2633 r0 *1 743.155,1129.05 rfnmoshv
2633$2633 \$1349 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2634 r0 *1 744.395,1129.05 rfnmoshv
2634$2634 IOVSS|VSS \$1145 \$1350 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2635 r0 *1 746.175,1129.05 rfnmoshv
2635$2635 \$1350 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2636 r0 *1 747.415,1129.05 rfnmoshv
2636$2636 IOVSS|VSS \$1145 \$1351 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2637 r0 *1 749.195,1129.05 rfnmoshv
2637$2637 \$1351 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2638 r0 *1 750.435,1129.05 rfnmoshv
2638$2638 IOVSS|VSS \$1145 \$1352 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2639 r0 *1 752.215,1129.05 rfnmoshv
2639$2639 \$1352 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2640 r0 *1 753.455,1129.05 rfnmoshv
2640$2640 IOVSS|VSS \$1145 \$1353 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2641 r0 *1 755.235,1129.05 rfnmoshv
2641$2641 \$1353 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2642 r0 *1 756.475,1129.05 rfnmoshv
2642$2642 IOVSS|VSS \$1145 \$1354 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2643 r0 *1 758.255,1129.05 rfnmoshv
2643$2643 \$1354 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2644 r0 *1 759.495,1129.05 rfnmoshv
2644$2644 IOVSS|VSS \$1145 \$1355 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2645 r0 *1 761.275,1129.05 rfnmoshv
2645$2645 \$1355 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2646 r0 *1 762.515,1129.05 rfnmoshv
2646$2646 IOVSS|VSS \$1145 \$1356 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2647 r0 *1 764.295,1129.05 rfnmoshv
2647$2647 \$1356 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2648 r0 *1 765.535,1129.05 rfnmoshv
2648$2648 IOVSS|VSS \$1145 \$1357 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2649 r0 *1 767.315,1129.05 rfnmoshv
2649$2649 \$1357 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2650 r0 *1 768.555,1129.05 rfnmoshv
2650$2650 IOVSS|VSS \$1145 \$1358 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2651 r0 *1 770.335,1129.05 rfnmoshv
2651$2651 \$1358 \$1145 IOVSS|VSS IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2652 r0 *1 771.575,1129.05 rfnmoshv
2652$2652 IOVSS|VSS \$1145 \$1359 IOVSS|VSS rfnmoshv W=4.3999999999999995
+ L=0.5999999999999998
* device instance $2653 r0 *1 865.09,598.44 rfpmoshv
2653$2653 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2654 r0 *1 865.09,599.32 rfpmoshv
2654$2654 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2655 r0 *1 865.09,600.2 rfpmoshv
2655$2655 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2656 r0 *1 865.09,601.08 rfpmoshv
2656$2656 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2657 r0 *1 865.09,601.96 rfpmoshv
2657$2657 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2658 r0 *1 865.09,602.84 rfpmoshv
2658$2658 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2659 r0 *1 865.09,603.72 rfpmoshv
2659$2659 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2660 r0 *1 865.09,604.6 rfpmoshv
2660$2660 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2661 r0 *1 865.09,605.48 rfpmoshv
2661$2661 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2662 r0 *1 865.09,606.36 rfpmoshv
2662$2662 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2663 r0 *1 865.09,607.24 rfpmoshv
2663$2663 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2664 r0 *1 865.09,608.12 rfpmoshv
2664$2664 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2665 r0 *1 865.09,609 rfpmoshv
2665$2665 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2666 r0 *1 865.09,609.88 rfpmoshv
2666$2666 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2667 r0 *1 865.09,610.76 rfpmoshv
2667$2667 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2668 r0 *1 865.09,611.64 rfpmoshv
2668$2668 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2669 r0 *1 865.09,612.52 rfpmoshv
2669$2669 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2670 r0 *1 865.09,613.4 rfpmoshv
2670$2670 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2671 r0 *1 865.09,614.28 rfpmoshv
2671$2671 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2672 r0 *1 865.09,615.16 rfpmoshv
2672$2672 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2673 r0 *1 865.09,616.04 rfpmoshv
2673$2673 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2674 r0 *1 865.09,616.92 rfpmoshv
2674$2674 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2675 r0 *1 865.09,617.8 rfpmoshv
2675$2675 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2676 r0 *1 865.09,618.68 rfpmoshv
2676$2676 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2677 r0 *1 865.09,619.56 rfpmoshv
2677$2677 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2678 r0 *1 865.09,620.44 rfpmoshv
2678$2678 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2679 r0 *1 865.09,621.32 rfpmoshv
2679$2679 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2680 r0 *1 865.09,622.2 rfpmoshv
2680$2680 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2681 r0 *1 865.09,623.08 rfpmoshv
2681$2681 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2682 r0 *1 865.09,623.96 rfpmoshv
2682$2682 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2683 r0 *1 865.09,624.84 rfpmoshv
2683$2683 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2684 r0 *1 865.09,625.72 rfpmoshv
2684$2684 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2685 r0 *1 865.09,626.6 rfpmoshv
2685$2685 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2686 r0 *1 865.09,627.48 rfpmoshv
2686$2686 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2687 r0 *1 865.09,628.36 rfpmoshv
2687$2687 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2688 r0 *1 865.09,629.24 rfpmoshv
2688$2688 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2689 r0 *1 865.09,630.12 rfpmoshv
2689$2689 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2690 r0 *1 865.09,631 rfpmoshv
2690$2690 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2691 r0 *1 865.09,631.88 rfpmoshv
2691$2691 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2692 r0 *1 865.09,632.76 rfpmoshv
2692$2692 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2693 r0 *1 865.09,633.64 rfpmoshv
2693$2693 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2694 r0 *1 865.09,634.52 rfpmoshv
2694$2694 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2695 r0 *1 865.09,635.4 rfpmoshv
2695$2695 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2696 r0 *1 865.09,636.28 rfpmoshv
2696$2696 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2697 r0 *1 865.09,637.16 rfpmoshv
2697$2697 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2698 r0 *1 865.09,638.04 rfpmoshv
2698$2698 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2699 r0 *1 865.09,638.92 rfpmoshv
2699$2699 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2700 r0 *1 865.09,639.8 rfpmoshv
2700$2700 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2701 r0 *1 865.09,640.68 rfpmoshv
2701$2701 IOVDD IOVDD \$626 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2702 r0 *1 865.09,641.56 rfpmoshv
2702$2702 \$626 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2703 r0 *1 18.44,1045.09 rfpmoshv
2703$2703 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2704 r0 *1 19.32,1045.09 rfpmoshv
2704$2704 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2705 r0 *1 20.2,1045.09 rfpmoshv
2705$2705 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2706 r0 *1 21.08,1045.09 rfpmoshv
2706$2706 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2707 r0 *1 21.96,1045.09 rfpmoshv
2707$2707 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2708 r0 *1 22.84,1045.09 rfpmoshv
2708$2708 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2709 r0 *1 23.72,1045.09 rfpmoshv
2709$2709 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2710 r0 *1 24.6,1045.09 rfpmoshv
2710$2710 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2711 r0 *1 25.48,1045.09 rfpmoshv
2711$2711 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2712 r0 *1 26.36,1045.09 rfpmoshv
2712$2712 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2713 r0 *1 27.24,1045.09 rfpmoshv
2713$2713 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2714 r0 *1 28.12,1045.09 rfpmoshv
2714$2714 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2715 r0 *1 29,1045.09 rfpmoshv
2715$2715 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2716 r0 *1 29.88,1045.09 rfpmoshv
2716$2716 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2717 r0 *1 30.76,1045.09 rfpmoshv
2717$2717 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2718 r0 *1 31.64,1045.09 rfpmoshv
2718$2718 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2719 r0 *1 32.52,1045.09 rfpmoshv
2719$2719 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2720 r0 *1 33.4,1045.09 rfpmoshv
2720$2720 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2721 r0 *1 34.28,1045.09 rfpmoshv
2721$2721 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2722 r0 *1 35.16,1045.09 rfpmoshv
2722$2722 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2723 r0 *1 36.04,1045.09 rfpmoshv
2723$2723 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2724 r0 *1 36.92,1045.09 rfpmoshv
2724$2724 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2725 r0 *1 37.8,1045.09 rfpmoshv
2725$2725 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2726 r0 *1 38.68,1045.09 rfpmoshv
2726$2726 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2727 r0 *1 39.56,1045.09 rfpmoshv
2727$2727 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2728 r0 *1 40.44,1045.09 rfpmoshv
2728$2728 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2729 r0 *1 41.32,1045.09 rfpmoshv
2729$2729 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2730 r0 *1 42.2,1045.09 rfpmoshv
2730$2730 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2731 r0 *1 43.08,1045.09 rfpmoshv
2731$2731 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2732 r0 *1 43.96,1045.09 rfpmoshv
2732$2732 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2733 r0 *1 44.84,1045.09 rfpmoshv
2733$2733 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2734 r0 *1 45.72,1045.09 rfpmoshv
2734$2734 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2735 r0 *1 46.6,1045.09 rfpmoshv
2735$2735 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2736 r0 *1 47.48,1045.09 rfpmoshv
2736$2736 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2737 r0 *1 48.36,1045.09 rfpmoshv
2737$2737 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2738 r0 *1 49.24,1045.09 rfpmoshv
2738$2738 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2739 r0 *1 50.12,1045.09 rfpmoshv
2739$2739 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2740 r0 *1 51,1045.09 rfpmoshv
2740$2740 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2741 r0 *1 51.88,1045.09 rfpmoshv
2741$2741 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2742 r0 *1 52.76,1045.09 rfpmoshv
2742$2742 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2743 r0 *1 53.64,1045.09 rfpmoshv
2743$2743 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2744 r0 *1 54.52,1045.09 rfpmoshv
2744$2744 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2745 r0 *1 55.4,1045.09 rfpmoshv
2745$2745 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2746 r0 *1 56.28,1045.09 rfpmoshv
2746$2746 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2747 r0 *1 57.16,1045.09 rfpmoshv
2747$2747 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2748 r0 *1 58.04,1045.09 rfpmoshv
2748$2748 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2749 r0 *1 58.92,1045.09 rfpmoshv
2749$2749 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2750 r0 *1 59.8,1045.09 rfpmoshv
2750$2750 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2751 r0 *1 60.68,1045.09 rfpmoshv
2751$2751 AVDD|IOVDD AVDD|IOVDD \$1143 AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2752 r0 *1 61.56,1045.09 rfpmoshv
2752$2752 \$1143 AVDD|IOVDD AVDD|IOVDD AVDD|IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2753 r0 *1 318.44,1045.09 rfpmoshv
2753$2753 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2754 r0 *1 319.32,1045.09 rfpmoshv
2754$2754 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2755 r0 *1 320.2,1045.09 rfpmoshv
2755$2755 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2756 r0 *1 321.08,1045.09 rfpmoshv
2756$2756 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2757 r0 *1 321.96,1045.09 rfpmoshv
2757$2757 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2758 r0 *1 322.84,1045.09 rfpmoshv
2758$2758 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2759 r0 *1 323.72,1045.09 rfpmoshv
2759$2759 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2760 r0 *1 324.6,1045.09 rfpmoshv
2760$2760 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2761 r0 *1 325.48,1045.09 rfpmoshv
2761$2761 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2762 r0 *1 326.36,1045.09 rfpmoshv
2762$2762 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2763 r0 *1 327.24,1045.09 rfpmoshv
2763$2763 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2764 r0 *1 328.12,1045.09 rfpmoshv
2764$2764 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2765 r0 *1 329,1045.09 rfpmoshv
2765$2765 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2766 r0 *1 329.88,1045.09 rfpmoshv
2766$2766 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2767 r0 *1 330.76,1045.09 rfpmoshv
2767$2767 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2768 r0 *1 331.64,1045.09 rfpmoshv
2768$2768 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2769 r0 *1 332.52,1045.09 rfpmoshv
2769$2769 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2770 r0 *1 333.4,1045.09 rfpmoshv
2770$2770 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2771 r0 *1 334.28,1045.09 rfpmoshv
2771$2771 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2772 r0 *1 335.16,1045.09 rfpmoshv
2772$2772 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2773 r0 *1 336.04,1045.09 rfpmoshv
2773$2773 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2774 r0 *1 336.92,1045.09 rfpmoshv
2774$2774 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2775 r0 *1 337.8,1045.09 rfpmoshv
2775$2775 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2776 r0 *1 338.68,1045.09 rfpmoshv
2776$2776 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2777 r0 *1 339.56,1045.09 rfpmoshv
2777$2777 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2778 r0 *1 340.44,1045.09 rfpmoshv
2778$2778 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2779 r0 *1 341.32,1045.09 rfpmoshv
2779$2779 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2780 r0 *1 342.2,1045.09 rfpmoshv
2780$2780 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2781 r0 *1 343.08,1045.09 rfpmoshv
2781$2781 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2782 r0 *1 343.96,1045.09 rfpmoshv
2782$2782 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2783 r0 *1 344.84,1045.09 rfpmoshv
2783$2783 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2784 r0 *1 345.72,1045.09 rfpmoshv
2784$2784 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2785 r0 *1 346.6,1045.09 rfpmoshv
2785$2785 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2786 r0 *1 347.48,1045.09 rfpmoshv
2786$2786 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2787 r0 *1 348.36,1045.09 rfpmoshv
2787$2787 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2788 r0 *1 349.24,1045.09 rfpmoshv
2788$2788 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2789 r0 *1 350.12,1045.09 rfpmoshv
2789$2789 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2790 r0 *1 351,1045.09 rfpmoshv
2790$2790 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2791 r0 *1 351.88,1045.09 rfpmoshv
2791$2791 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2792 r0 *1 352.76,1045.09 rfpmoshv
2792$2792 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2793 r0 *1 353.64,1045.09 rfpmoshv
2793$2793 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2794 r0 *1 354.52,1045.09 rfpmoshv
2794$2794 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2795 r0 *1 355.4,1045.09 rfpmoshv
2795$2795 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2796 r0 *1 356.28,1045.09 rfpmoshv
2796$2796 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2797 r0 *1 357.16,1045.09 rfpmoshv
2797$2797 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2798 r0 *1 358.04,1045.09 rfpmoshv
2798$2798 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2799 r0 *1 358.92,1045.09 rfpmoshv
2799$2799 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2800 r0 *1 359.8,1045.09 rfpmoshv
2800$2800 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2801 r0 *1 360.68,1045.09 rfpmoshv
2801$2801 IOVDD IOVDD \$1144 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2802 r0 *1 361.56,1045.09 rfpmoshv
2802$2802 \$1144 IOVDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2803 r0 *1 718.44,1045.09 rfpmoshv
2803$2803 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2804 r0 *1 719.32,1045.09 rfpmoshv
2804$2804 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2805 r0 *1 720.2,1045.09 rfpmoshv
2805$2805 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2806 r0 *1 721.08,1045.09 rfpmoshv
2806$2806 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2807 r0 *1 721.96,1045.09 rfpmoshv
2807$2807 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2808 r0 *1 722.84,1045.09 rfpmoshv
2808$2808 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2809 r0 *1 723.72,1045.09 rfpmoshv
2809$2809 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2810 r0 *1 724.6,1045.09 rfpmoshv
2810$2810 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2811 r0 *1 725.48,1045.09 rfpmoshv
2811$2811 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2812 r0 *1 726.36,1045.09 rfpmoshv
2812$2812 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2813 r0 *1 727.24,1045.09 rfpmoshv
2813$2813 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2814 r0 *1 728.12,1045.09 rfpmoshv
2814$2814 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2815 r0 *1 729,1045.09 rfpmoshv
2815$2815 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2816 r0 *1 729.88,1045.09 rfpmoshv
2816$2816 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2817 r0 *1 730.76,1045.09 rfpmoshv
2817$2817 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2818 r0 *1 731.64,1045.09 rfpmoshv
2818$2818 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2819 r0 *1 732.52,1045.09 rfpmoshv
2819$2819 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2820 r0 *1 733.4,1045.09 rfpmoshv
2820$2820 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2821 r0 *1 734.28,1045.09 rfpmoshv
2821$2821 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2822 r0 *1 735.16,1045.09 rfpmoshv
2822$2822 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2823 r0 *1 736.04,1045.09 rfpmoshv
2823$2823 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2824 r0 *1 736.92,1045.09 rfpmoshv
2824$2824 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2825 r0 *1 737.8,1045.09 rfpmoshv
2825$2825 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2826 r0 *1 738.68,1045.09 rfpmoshv
2826$2826 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2827 r0 *1 739.56,1045.09 rfpmoshv
2827$2827 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2828 r0 *1 740.44,1045.09 rfpmoshv
2828$2828 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2829 r0 *1 741.32,1045.09 rfpmoshv
2829$2829 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2830 r0 *1 742.2,1045.09 rfpmoshv
2830$2830 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2831 r0 *1 743.08,1045.09 rfpmoshv
2831$2831 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2832 r0 *1 743.96,1045.09 rfpmoshv
2832$2832 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2833 r0 *1 744.84,1045.09 rfpmoshv
2833$2833 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2834 r0 *1 745.72,1045.09 rfpmoshv
2834$2834 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2835 r0 *1 746.6,1045.09 rfpmoshv
2835$2835 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2836 r0 *1 747.48,1045.09 rfpmoshv
2836$2836 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2837 r0 *1 748.36,1045.09 rfpmoshv
2837$2837 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2838 r0 *1 749.24,1045.09 rfpmoshv
2838$2838 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2839 r0 *1 750.12,1045.09 rfpmoshv
2839$2839 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2840 r0 *1 751,1045.09 rfpmoshv
2840$2840 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2841 r0 *1 751.88,1045.09 rfpmoshv
2841$2841 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2842 r0 *1 752.76,1045.09 rfpmoshv
2842$2842 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2843 r0 *1 753.64,1045.09 rfpmoshv
2843$2843 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2844 r0 *1 754.52,1045.09 rfpmoshv
2844$2844 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2845 r0 *1 755.4,1045.09 rfpmoshv
2845$2845 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2846 r0 *1 756.28,1045.09 rfpmoshv
2846$2846 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2847 r0 *1 757.16,1045.09 rfpmoshv
2847$2847 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2848 r0 *1 758.04,1045.09 rfpmoshv
2848$2848 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2849 r0 *1 758.92,1045.09 rfpmoshv
2849$2849 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2850 r0 *1 759.8,1045.09 rfpmoshv
2850$2850 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2851 r0 *1 760.68,1045.09 rfpmoshv
2851$2851 IOVDD VDD \$1145 IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2852 r0 *1 761.56,1045.09 rfpmoshv
2852$2852 \$1145 VDD IOVDD IOVDD rfpmoshv W=6.999999999999998
+ L=0.4999999999999999
* device instance $2853 r0 *1 4.54,24.19 dantenna
D$2853 IOVSS|VSS IOVSS|VSS dantenna A=35.0028 P=58.08 m=1
* device instance $2854 r0 *1 9.04,24.19 dantenna
D$2854 IOVSS|VSS IOVSS|VSS dantenna A=35.0028 P=58.08 m=1
* device instance $2855 r0 *1 104.54,24.19 dantenna
D$2855 IOVSS|VSS IOVSS|VSS dantenna A=35.0028 P=58.08 m=1
* device instance $2856 r0 *1 109.04,24.19 dantenna
D$2856 IOVSS|VSS IOVSS|VSS dantenna A=35.0028 P=58.08 m=1
* device instance $2857 r0 *1 204.54,24.19 dantenna
D$2857 IOVSS|VSS RES dantenna A=35.0028 P=58.08 m=1
* device instance $2858 r0 *1 209.04,24.19 dantenna
D$2858 IOVSS|VSS RES dantenna A=35.0028 P=58.08 m=1
* device instance $2859 r0 *1 304.54,24.19 dantenna
D$2859 IOVSS|VSS IOVSS|VSS dantenna A=35.0028 P=58.08 m=1
* device instance $2860 r0 *1 309.04,24.19 dantenna
D$2860 IOVSS|VSS IOVSS|VSS dantenna A=35.0028 P=58.08 m=1
* device instance $2861 r0 *1 404.54,24.19 dantenna
D$2861 IOVSS|VSS CK4 dantenna A=35.0028 P=58.08 m=1
* device instance $2862 r0 *1 409.04,24.19 dantenna
D$2862 IOVSS|VSS CK4 dantenna A=35.0028 P=58.08 m=1
* device instance $2863 r0 *1 504.54,24.19 dantenna
D$2863 IOVSS|VSS CK5 dantenna A=35.0028 P=58.08 m=1
* device instance $2864 r0 *1 509.04,24.19 dantenna
D$2864 IOVSS|VSS CK5 dantenna A=35.0028 P=58.08 m=1
* device instance $2865 r0 *1 604.54,24.19 dantenna
D$2865 IOVSS|VSS CK6 dantenna A=35.0028 P=58.08 m=1
* device instance $2866 r0 *1 609.04,24.19 dantenna
D$2866 IOVSS|VSS CK6 dantenna A=35.0028 P=58.08 m=1
* device instance $2867 r0 *1 704.54,24.19 dantenna
D$2867 IOVSS|VSS IOVSS|VSS dantenna A=35.0028 P=58.08 m=1
* device instance $2868 r0 *1 709.04,24.19 dantenna
D$2868 IOVSS|VSS IOVSS|VSS dantenna A=35.0028 P=58.08 m=1
* device instance $2869 r0 *1 -159.56,320 dantenna
D$2869 IOVSS|VSS IN5|PAD dantenna A=35.0028 P=58.08 m=1
* device instance $2870 r0 *1 -159.56,220 dantenna
D$2870 IOVSS|VSS IN6|PAD dantenna A=35.0028 P=58.08 m=1
* device instance $2871 r0 *1 -155.06,320 dantenna
D$2871 IOVSS|VSS IN5|PAD dantenna A=35.0028 P=58.08 m=1
* device instance $2872 r0 *1 -155.06,220 dantenna
D$2872 IOVSS|VSS IN6|PAD dantenna A=35.0028 P=58.08 m=1
* device instance $2873 r0 *1 -37.46,337.63 dantenna
D$2873 IOVSS|VSS PADRES|in5_c dantenna A=1.984 P=7.48 m=1
* device instance $2874 r0 *1 -37.46,237.63 dantenna
D$2874 IOVSS|VSS PADRES|in6_c dantenna A=1.984 P=7.48 m=1
* device instance $2875 r0 *1 245.225,142.54 dantenna
D$2875 IOVSS|VSS \$129 dantenna A=1.984 P=7.48 m=1
* device instance $2876 r0 *1 445.225,142.54 dantenna
D$2876 IOVSS|VSS \$130 dantenna A=1.984 P=7.48 m=1
* device instance $2877 r0 *1 545.225,142.54 dantenna
D$2877 IOVSS|VSS \$132 dantenna A=1.984 P=7.48 m=1
* device instance $2878 r0 *1 645.225,142.54 dantenna
D$2878 IOVSS|VSS \$133 dantenna A=1.984 P=7.48 m=1
* device instance $2879 r0 *1 935.06,220 dantenna
D$2879 IOVSS|VSS OUT6 dantenna A=35.0028 P=58.08 m=1
* device instance $2880 r0 *1 935.06,320 dantenna
D$2880 IOVSS|VSS OUT5 dantenna A=35.0028 P=58.08 m=1
* device instance $2881 r0 *1 939.56,320 dantenna
D$2881 IOVSS|VSS OUT5 dantenna A=35.0028 P=58.08 m=1
* device instance $2882 r0 *1 939.56,220 dantenna
D$2882 IOVSS|VSS OUT6 dantenna A=35.0028 P=58.08 m=1
* device instance $2883 r0 *1 947.17,297.975 dantenna
D$2883 IOVSS|VSS \$366 dantenna A=0.192 P=1.88 m=1
* device instance $2884 r0 *1 947.17,197.975 dantenna
D$2884 IOVSS|VSS \$253 dantenna A=0.192 P=1.88 m=1
* device instance $2885 r0 *1 947.17,397.975 dantenna
D$2885 IOVSS|VSS \$479 dantenna A=0.192 P=1.88 m=1
* device instance $2886 r0 *1 -159.56,420 dantenna
D$2886 IOVSS|VSS IN4|PAD dantenna A=35.0028 P=58.08 m=1
* device instance $2887 r0 *1 -155.06,420 dantenna
D$2887 IOVSS|VSS IN4|PAD dantenna A=35.0028 P=58.08 m=1
* device instance $2888 r0 *1 935.06,420 dantenna
D$2888 IOVSS|VSS OUT4 dantenna A=35.0028 P=58.08 m=1
* device instance $2889 r0 *1 939.56,420 dantenna
D$2889 IOVSS|VSS OUT4 dantenna A=35.0028 P=58.08 m=1
* device instance $2890 r0 *1 -37.46,437.63 dantenna
D$2890 IOVSS|VSS PADRES|in4_c dantenna A=1.984 P=7.48 m=1
* device instance $2891 r0 *1 935.81,484.54 dantenna
D$2891 IOVSS|VSS IOVSS|VSS dantenna A=35.0028 P=58.08 m=1
* device instance $2892 r0 *1 935.81,489.04 dantenna
D$2892 IOVSS|VSS IOVSS|VSS dantenna A=35.0028 P=58.08 m=1
* device instance $2893 r0 *1 -159.56,520 dantenna
D$2893 IOVSS|VSS PAD|VLO dantenna A=35.0028 P=58.08 m=1
* device instance $2894 r0 *1 -155.06,520 dantenna
D$2894 IOVSS|VSS PAD|VLO dantenna A=35.0028 P=58.08 m=1
* device instance $2895 r0 *1 -37.46,537.63 dantenna
D$2895 IOVSS|VSS PADRES dantenna A=1.984 P=7.48 m=1
* device instance $2896 r0 *1 932.65,584.765 dantenna
D$2896 IOVSS|VSS \$626 dantenna A=0.192 P=1.88 m=1
* device instance $2897 r0 *1 -159.56,620 dantenna
D$2897 IOVSS|VSS PAD|VHI dantenna A=35.0028 P=58.08 m=1
* device instance $2898 r0 *1 -155.06,620 dantenna
D$2898 IOVSS|VSS PAD|VHI dantenna A=35.0028 P=58.08 m=1
* device instance $2899 r0 *1 -37.46,637.63 dantenna
D$2899 IOVSS|VSS PADRES$1 dantenna A=1.984 P=7.48 m=1
* device instance $2900 r0 *1 947.17,697.975 dantenna
D$2900 IOVSS|VSS \$766 dantenna A=0.192 P=1.88 m=1
* device instance $2901 r0 *1 -159.56,720 dantenna
D$2901 IOVSS|VSS IN3|PAD dantenna A=35.0028 P=58.08 m=1
* device instance $2902 r0 *1 -155.06,720 dantenna
D$2902 IOVSS|VSS IN3|PAD dantenna A=35.0028 P=58.08 m=1
* device instance $2903 r0 *1 935.06,720 dantenna
D$2903 IOVSS|VSS OUT3 dantenna A=35.0028 P=58.08 m=1
* device instance $2904 r0 *1 939.56,720 dantenna
D$2904 IOVSS|VSS OUT3 dantenna A=35.0028 P=58.08 m=1
* device instance $2905 r0 *1 -37.46,737.63 dantenna
D$2905 IOVSS|VSS PADRES|in3_c dantenna A=1.984 P=7.48 m=1
* device instance $2906 r0 *1 947.17,797.975 dantenna
D$2906 IOVSS|VSS \$879 dantenna A=0.192 P=1.88 m=1
* device instance $2907 r0 *1 -159.56,820 dantenna
D$2907 IOVSS|VSS IN2|PAD dantenna A=35.0028 P=58.08 m=1
* device instance $2908 r0 *1 -155.06,820 dantenna
D$2908 IOVSS|VSS IN2|PAD dantenna A=35.0028 P=58.08 m=1
* device instance $2909 r0 *1 935.06,820 dantenna
D$2909 IOVSS|VSS OUT2 dantenna A=35.0028 P=58.08 m=1
* device instance $2910 r0 *1 939.56,820 dantenna
D$2910 IOVSS|VSS OUT2 dantenna A=35.0028 P=58.08 m=1
* device instance $2911 r0 *1 -37.46,837.63 dantenna
D$2911 IOVSS|VSS PADRES|in2_c dantenna A=1.984 P=7.48 m=1
* device instance $2912 r0 *1 947.17,897.975 dantenna
D$2912 IOVSS|VSS \$992 dantenna A=0.192 P=1.88 m=1
* device instance $2913 r0 *1 -159.56,920 dantenna
D$2913 IOVSS|VSS IN1|PAD dantenna A=35.0028 P=58.08 m=1
* device instance $2914 r0 *1 -155.06,920 dantenna
D$2914 IOVSS|VSS IN1|PAD dantenna A=35.0028 P=58.08 m=1
* device instance $2915 r0 *1 935.06,920 dantenna
D$2915 IOVSS|VSS OUT1 dantenna A=35.0028 P=58.08 m=1
* device instance $2916 r0 *1 939.56,920 dantenna
D$2916 IOVSS|VSS OUT1 dantenna A=35.0028 P=58.08 m=1
* device instance $2917 r0 *1 -37.46,937.63 dantenna
D$2917 IOVSS|VSS PADRES|in1_c dantenna A=1.984 P=7.48 m=1
* device instance $2918 r0 *1 157.63,997.46 dantenna
D$2918 IOVSS|VSS PADRES|vref_c dantenna A=1.984 P=7.48 m=1
* device instance $2919 r0 *1 257.63,997.46 dantenna
D$2919 IOVSS|VSS PADRES$2 dantenna A=1.984 P=7.48 m=1
* device instance $2920 r0 *1 445.225,997.46 dantenna
D$2920 IOVSS|VSS \$1070 dantenna A=1.984 P=7.48 m=1
* device instance $2921 r0 *1 545.225,997.46 dantenna
D$2921 IOVSS|VSS \$1071 dantenna A=1.984 P=7.48 m=1
* device instance $2922 r0 *1 645.225,997.46 dantenna
D$2922 IOVSS|VSS \$1072 dantenna A=1.984 P=7.48 m=1
* device instance $2923 r0 *1 404.54,1115.81 dantenna
D$2923 IOVSS|VSS CK3 dantenna A=35.0028 P=58.08 m=1
* device instance $2924 r0 *1 409.04,1115.81 dantenna
D$2924 IOVSS|VSS CK3 dantenna A=35.0028 P=58.08 m=1
* device instance $2925 r0 *1 504.54,1115.81 dantenna
D$2925 IOVSS|VSS CK2 dantenna A=35.0028 P=58.08 m=1
* device instance $2926 r0 *1 509.04,1115.81 dantenna
D$2926 IOVSS|VSS CK2 dantenna A=35.0028 P=58.08 m=1
* device instance $2927 r0 *1 604.54,1115.81 dantenna
D$2927 IOVSS|VSS CK1 dantenna A=35.0028 P=58.08 m=1
* device instance $2928 r0 *1 609.04,1115.81 dantenna
D$2928 IOVSS|VSS CK1 dantenna A=35.0028 P=58.08 m=1
* device instance $2929 r0 *1 4.765,1112.65 dantenna
D$2929 IOVSS|VSS \$1143 dantenna A=0.192 P=1.88 m=1
* device instance $2930 r0 *1 140,1115.06 dantenna
D$2930 IOVSS|VSS PAD|VREF dantenna A=35.0028 P=58.08 m=1
* device instance $2931 r0 *1 240,1115.06 dantenna
D$2931 IOVSS|VSS PAD|VLDO dantenna A=35.0028 P=58.08 m=1
* device instance $2932 r0 *1 304.765,1112.65 dantenna
D$2932 IOVSS|VSS \$1144 dantenna A=0.192 P=1.88 m=1
* device instance $2933 r0 *1 704.765,1112.65 dantenna
D$2933 IOVSS|VSS \$1145 dantenna A=0.192 P=1.88 m=1
* device instance $2934 r0 *1 140,1119.56 dantenna
D$2934 IOVSS|VSS PAD|VREF dantenna A=35.0028 P=58.08 m=1
* device instance $2935 r0 *1 240,1119.56 dantenna
D$2935 IOVSS|VSS PAD|VLDO dantenna A=35.0028 P=58.08 m=1
* device instance $2936 r0 *1 4.54,83.19 dpantenna
D$2936 IOVSS|VSS AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2937 r0 *1 9.04,83.19 dpantenna
D$2937 IOVSS|VSS AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2938 r0 *1 104.54,83.19 dpantenna
D$2938 IOVSS|VSS AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2939 r0 *1 109.04,83.19 dpantenna
D$2939 IOVSS|VSS AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2940 r0 *1 204.54,83.19 dpantenna
D$2940 RES IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2941 r0 *1 209.04,83.19 dpantenna
D$2941 RES IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2942 r0 *1 304.54,83.19 dpantenna
D$2942 IOVSS|VSS IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2943 r0 *1 309.04,83.19 dpantenna
D$2943 IOVSS|VSS IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2944 r0 *1 404.54,83.19 dpantenna
D$2944 CK4 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2945 r0 *1 409.04,83.19 dpantenna
D$2945 CK4 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2946 r0 *1 504.54,83.19 dpantenna
D$2946 CK5 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2947 r0 *1 509.04,83.19 dpantenna
D$2947 CK5 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2948 r0 *1 604.54,83.19 dpantenna
D$2948 CK6 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2949 r0 *1 609.04,83.19 dpantenna
D$2949 CK6 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2950 r0 *1 704.54,83.19 dpantenna
D$2950 IOVSS|VSS IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2951 r0 *1 709.04,83.19 dpantenna
D$2951 IOVSS|VSS IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2952 r0 *1 -124.04,320 dpantenna
D$2952 IN5|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2953 r0 *1 -124.04,220 dpantenna
D$2953 IN6|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2954 r0 *1 -119.54,320 dpantenna
D$2954 IN5|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2955 r0 *1 -119.54,220 dpantenna
D$2955 IN6|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2956 r0 *1 -32.49,335.46 dpantenna
D$2956 PADRES|in5_c AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2957 r0 *1 -32.49,235.46 dpantenna
D$2957 PADRES|in6_c AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2958 r0 *1 243.055,147.51 dpantenna
D$2958 \$129 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2959 r0 *1 443.055,147.51 dpantenna
D$2959 \$130 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2960 r0 *1 543.055,147.51 dpantenna
D$2960 \$132 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2961 r0 *1 643.055,147.51 dpantenna
D$2961 \$133 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2962 r0 *1 878.81,197.975 dpantenna
D$2962 \$218 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $2963 r0 *1 878.81,297.975 dpantenna
D$2963 \$331 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $2964 r0 *1 899.54,320 dpantenna
D$2964 OUT5 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2965 r0 *1 899.54,220 dpantenna
D$2965 OUT6 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2966 r0 *1 904.04,220 dpantenna
D$2966 OUT6 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2967 r0 *1 904.04,320 dpantenna
D$2967 OUT5 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2968 r0 *1 -124.04,420 dpantenna
D$2968 IN4|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2969 r0 *1 -119.54,420 dpantenna
D$2969 IN4|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2970 r0 *1 878.81,397.975 dpantenna
D$2970 \$444 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $2971 r0 *1 899.54,420 dpantenna
D$2971 OUT4 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2972 r0 *1 904.04,420 dpantenna
D$2972 OUT4 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2973 r0 *1 -32.49,435.46 dpantenna
D$2973 PADRES|in4_c AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2974 r0 *1 876.81,484.54 dpantenna
D$2974 IOVSS|VSS IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2975 r0 *1 876.81,489.04 dpantenna
D$2975 IOVSS|VSS IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2976 r0 *1 -124.04,520 dpantenna
D$2976 PAD|VLO AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2977 r0 *1 -119.54,520 dpantenna
D$2977 PAD|VLO AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2978 r0 *1 -32.49,535.46 dpantenna
D$2978 PADRES AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2979 r0 *1 -124.04,620 dpantenna
D$2979 PAD|VHI AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2980 r0 *1 -119.54,620 dpantenna
D$2980 PAD|VHI AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2981 r0 *1 -32.49,635.46 dpantenna
D$2981 PADRES$1 AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2982 r0 *1 878.81,697.975 dpantenna
D$2982 \$731 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $2983 r0 *1 -124.04,720 dpantenna
D$2983 IN3|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2984 r0 *1 -119.54,720 dpantenna
D$2984 IN3|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2985 r0 *1 899.54,720 dpantenna
D$2985 OUT3 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2986 r0 *1 904.04,720 dpantenna
D$2986 OUT3 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2987 r0 *1 -32.49,735.46 dpantenna
D$2987 PADRES|in3_c AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2988 r0 *1 878.81,797.975 dpantenna
D$2988 \$844 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $2989 r0 *1 -124.04,820 dpantenna
D$2989 IN2|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2990 r0 *1 -119.54,820 dpantenna
D$2990 IN2|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2991 r0 *1 899.54,820 dpantenna
D$2991 OUT2 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2992 r0 *1 904.04,820 dpantenna
D$2992 OUT2 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2993 r0 *1 -32.49,835.46 dpantenna
D$2993 PADRES|in2_c AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2994 r0 *1 878.81,897.975 dpantenna
D$2994 \$957 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $2995 r0 *1 -124.04,920 dpantenna
D$2995 IN1|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2996 r0 *1 -119.54,920 dpantenna
D$2996 IN1|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2997 r0 *1 899.54,920 dpantenna
D$2997 OUT1 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2998 r0 *1 904.04,920 dpantenna
D$2998 OUT1 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $2999 r0 *1 -32.49,935.46 dpantenna
D$2999 PADRES|in1_c AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3000 r0 *1 155.46,992.49 dpantenna
D$3000 PADRES|vref_c AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3001 r0 *1 255.46,992.49 dpantenna
D$3001 PADRES$2 AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3002 r0 *1 443.055,992.49 dpantenna
D$3002 \$1070 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3003 r0 *1 543.055,992.49 dpantenna
D$3003 \$1071 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3004 r0 *1 643.055,992.49 dpantenna
D$3004 \$1072 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3005 r0 *1 404.54,1056.81 dpantenna
D$3005 CK3 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $3006 r0 *1 409.04,1056.81 dpantenna
D$3006 CK3 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $3007 r0 *1 504.54,1056.81 dpantenna
D$3007 CK2 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $3008 r0 *1 509.04,1056.81 dpantenna
D$3008 CK2 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $3009 r0 *1 604.54,1056.81 dpantenna
D$3009 CK1 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $3010 r0 *1 609.04,1056.81 dpantenna
D$3010 CK1 IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $3011 r0 *1 140,1084.04 dpantenna
D$3011 PAD|VREF AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $3012 r0 *1 140,1079.54 dpantenna
D$3012 PAD|VREF AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $3013 r0 *1 240,1084.04 dpantenna
D$3013 PAD|VLDO AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $3014 r0 *1 240,1079.54 dpantenna
D$3014 PAD|VLDO AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=1
* device instance $3015 r0 *1 240.685,141.11 res_rppd
R$3015 RES \$129 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $3016 r0 *1 440.685,141.11 res_rppd
R$3016 CK4 \$130 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $3017 r0 *1 540.685,141.11 res_rppd
R$3017 CK5 \$132 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $3018 r0 *1 640.685,141.11 res_rppd
R$3018 CK6 \$133 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $3019 r0 *1 -171.25,246.305 res_rppd
R$3019 IOVSS|VSS \$227 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $3020 r0 *1 -112.25,246.305 res_rppd
R$3020 AVDD|IOVDD \$228 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $3021 r0 *1 -38.89,233.09 res_rppd
R$3021 IN6|PAD PADRES|in6_c res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $3022 r0 *1 -171.25,346.305 res_rppd
R$3022 IOVSS|VSS \$340 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $3023 r0 *1 -112.25,346.305 res_rppd
R$3023 AVDD|IOVDD \$341 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $3024 r0 *1 -38.89,333.09 res_rppd
R$3024 IN5|PAD PADRES|in5_c res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $3025 r0 *1 -171.25,446.305 res_rppd
R$3025 IOVSS|VSS \$453 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $3026 r0 *1 -112.25,446.305 res_rppd
R$3026 AVDD|IOVDD \$454 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $3027 r0 *1 -38.89,433.09 res_rppd
R$3027 IN4|PAD PADRES|in4_c res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $3028 r0 *1 -171.25,546.305 res_rppd
R$3028 IOVSS|VSS \$568 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $3029 r0 *1 -112.25,546.305 res_rppd
R$3029 AVDD|IOVDD \$569 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $3030 r0 *1 -38.89,533.09 res_rppd
R$3030 PAD|VLO PADRES res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $3031 r0 *1 -171.25,646.305 res_rppd
R$3031 IOVSS|VSS \$638 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $3032 r0 *1 -112.25,646.305 res_rppd
R$3032 AVDD|IOVDD \$639 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $3033 r0 *1 -38.89,633.09 res_rppd
R$3033 PAD|VHI PADRES$1 res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $3034 r0 *1 -171.25,746.305 res_rppd
R$3034 IOVSS|VSS \$740 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $3035 r0 *1 -112.25,746.305 res_rppd
R$3035 AVDD|IOVDD \$741 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $3036 r0 *1 -38.89,733.09 res_rppd
R$3036 IN3|PAD PADRES|in3_c res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $3037 r0 *1 -171.25,846.305 res_rppd
R$3037 IOVSS|VSS \$853 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $3038 r0 *1 -112.25,846.305 res_rppd
R$3038 AVDD|IOVDD \$854 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $3039 r0 *1 -38.89,833.09 res_rppd
R$3039 IN2|PAD PADRES|in2_c res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $3040 r0 *1 -171.25,946.305 res_rppd
R$3040 IOVSS|VSS \$966 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $3041 r0 *1 -112.25,946.305 res_rppd
R$3041 AVDD|IOVDD \$967 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $3042 r0 *1 -38.89,933.09 res_rppd
R$3042 IN1|PAD PADRES|in1_c res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $3043 r0 *1 153.09,996.03 res_rppd
R$3043 PADRES|vref_c PAD|VREF res_rppd w=0.9999999999999998
+ l=1.9999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $3044 r0 *1 253.09,996.03 res_rppd
R$3044 PADRES$2 PAD|VLDO res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $3045 r0 *1 440.685,996.03 res_rppd
R$3045 \$1070 CK3 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $3046 r0 *1 540.685,996.03 res_rppd
R$3046 \$1071 CK2 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $3047 r0 *1 640.685,996.03 res_rppd
R$3047 \$1072 CK1 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $3048 r0 *1 166.305,1126.85 res_rppd
R$3048 \$1397 IOVSS|VSS res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $3049 r0 *1 166.305,1058.49 res_rppd
R$3049 \$1160 AVDD|IOVDD res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $3050 r0 *1 266.305,1126.85 res_rppd
R$3050 \$1398 IOVSS|VSS res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $3051 r0 *1 266.305,1058.49 res_rppd
R$3051 \$1161 AVDD|IOVDD res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
.ENDS padring

* Extracted by KLayout with SG13G2 LVS runset on : 06/05/2024 02:34

* cell integ_5_split2
* pin sub!
.SUBCKT integ_5_split2 sub!
* device instance $1 r0 *1 -2.782,-5.221 sg13_lv_nmos
M$1 \$5 \$3 \$9 sub! sg13_lv_nmos W=0.64 L=0.13
* device instance $2 r0 *1 -2.272,-5.221 sg13_lv_nmos
M$2 sub! \$7 \$9 sub! sg13_lv_nmos W=0.64 L=0.13
* device instance $3 r0 *1 -1.762,-5.271 sg13_lv_nmos
M$3 sub! \$5 \$6 sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $4 r0 *1 2.984,-4.327 sg13_lv_nmos
M$4 \$1 \$6 \$20 sub! sg13_lv_nmos W=0.5 L=0.13
* device instance $5 r0 *1 4.141,0.398 sg13_lv_nmos
M$5 \$21 \$17 \$20 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $6 r0 *1 -2.782,-3.581 sg13_lv_pmos
M$6 \$10 \$3 \$5 \$10 sg13_lv_pmos W=0.84 L=0.13
* device instance $7 r0 *1 -2.272,-3.581 sg13_lv_pmos
M$7 \$10 \$7 \$5 \$10 sg13_lv_pmos W=0.84 L=0.13
* device instance $8 r0 *1 -1.762,-3.721 sg13_lv_pmos
M$8 \$10 \$5 \$6 \$10 sg13_lv_pmos W=1.12 L=0.13
* device instance $9 r0 *1 -3.021,0.4 sg13_lv_pmos
M$9 \$20 \$19 \$21 \$13 sg13_lv_pmos W=6.0 L=0.12999999999999998
.ENDS integ_5_split2

* Extracted by KLayout with SG13G2 LVS runset on : 03/05/2024 20:27

* cell sg13g2_IOPadOut16mA
* pin sub!
.SUBCKT sg13g2_IOPadOut16mA sub!
* device instance $1 r0 *1 37.48,159.005 sg13_lv_nmos
M$1 \$44 \$45 sub! sub! sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $2 r0 *1 40.99,159.005 sg13_lv_nmos
M$2 \$46 \$45 sub! sub! sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $3 r0 *1 34.58,10.95 sg13_hv_nmos
M$3 sub! \$6 \$1 sub! sg13_hv_nmos W=35.199999999999996 L=0.5999999999999998
* device instance $11 r0 *1 37.64,155.32 sg13_hv_nmos
M$11 \$38 \$45 sub! sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $12 r0 *1 38.47,155.32 sg13_hv_nmos
M$12 sub! \$44 \$39 sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $13 r0 *1 39.81,155.32 sg13_hv_nmos
M$13 sub! \$39 \$6 sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $14 r0 *1 41.15,155.32 sg13_hv_nmos
M$14 \$40 \$45 sub! sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $15 r0 *1 41.98,155.32 sg13_hv_nmos
M$15 sub! \$46 \$41 sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $16 r0 *1 43.32,155.32 sg13_hv_nmos
M$16 sub! \$41 \$32 sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $17 r0 *1 37.48,163.995 sg13_lv_pmos
M$17 \$44 \$45 \$36 \$36 sg13_lv_pmos W=4.749999999999999 L=0.12999999999999998
* device instance $18 r0 *1 40.99,163.995 sg13_lv_pmos
M$18 \$46 \$45 \$36 \$36 sg13_lv_pmos W=4.749999999999999 L=0.12999999999999998
* device instance $19 r0 *1 34.58,71.08 sg13_hv_pmos
M$19 \$21 \$32 \$1 \$21 sg13_hv_pmos W=106.55999999999996 L=0.5999999999999999
* device instance $35 r0 *1 37.64,151.18 sg13_hv_pmos
M$35 \$38 \$39 \$21 \$21 sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $36 r0 *1 38.47,151.18 sg13_hv_pmos
M$36 \$21 \$38 \$39 \$21 sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $37 r0 *1 41.15,151.18 sg13_hv_pmos
M$37 \$40 \$41 \$21 \$21 sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $38 r0 *1 41.98,151.18 sg13_hv_pmos
M$38 \$21 \$40 \$41 \$21 sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $39 r0 *1 39.81,151.18 sg13_hv_pmos
M$39 \$21 \$39 \$6 \$21 sg13_hv_pmos W=3.899999999999999 L=0.4499999999999999
* device instance $40 r0 *1 43.32,151.18 sg13_hv_pmos
M$40 \$21 \$41 \$32 \$21 sg13_hv_pmos W=3.899999999999999 L=0.4499999999999999
* device instance $41 r0 *1 17.975,12.83 dantenna
D$41 sub! \$6 dantenna A=0.192 P=1.88 m=1
* device instance $42 r0 *1 40,20.44 dantenna
D$42 sub! \$1 dantenna A=35.0028 P=58.08 m=2
* device instance $44 r0 *1 40,55.96 dpantenna
D$44 \$1 \$21 dpantenna A=35.0028 P=58.08 m=2
* device instance $46 r0 *1 17.975,81.19 dpantenna
D$46 \$32 \$21 dpantenna A=0.192 P=1.88 m=1
.ENDS sg13g2_IOPadOut16mA

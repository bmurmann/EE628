* Extracted by KLayout with SG13G2 LVS runset on : 03/05/2024 20:17

* cell sg13g2_IOPadIn
* pin PAD
* pin CORE
* pin sub!
.SUBCKT sg13g2_IOPadIn PAD CORE sub!
* device instance $1 r0 *1 40.255,159.005 sg13_lv_nmos
M$1 \$35 \$37 sub! sub! sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $2 r0 *1 41.765,159.055 sg13_hv_nmos
M$2 sub! CORE \$37 sub! sg13_hv_nmos W=2.6499999999999995 L=0.4499999999999999
* device instance $3 r0 *1 40.255,163.995 sg13_lv_pmos
M$3 \$35 \$37 \$22 \$22 sg13_lv_pmos W=4.749999999999999 L=0.12999999999999998
* device instance $4 r0 *1 41.765,163.945 sg13_hv_pmos
M$4 \$22 CORE \$37 \$22 sg13_hv_pmos W=4.6499999999999995 L=0.44999999999999984
* device instance $5 r0 *1 4.54,24.19 dantenna
D$5 sub! PAD dantenna A=35.0028 P=58.08 m=2
* device instance $7 r0 *1 45.225,142.54 dantenna
D$7 sub! CORE dantenna A=1.984 P=7.48 m=1
* device instance $8 r0 *1 4.54,83.19 dpantenna
D$8 PAD \$15 dpantenna A=35.0028 P=58.08 m=2
* device instance $10 r0 *1 43.055,147.51 dpantenna
D$10 CORE \$15 dpantenna A=3.1872 P=11.24 m=1
* device instance $11 r0 *1 40.685,141.11 rppd
R$11 PAD CORE rppd w=1 l=2 ps=0 b=0 m=1
.ENDS sg13g2_IOPadIn

* Extracted by KLayout with SG13G2 LVS runset on : 03/05/2024 04:26

* cell sg13g2_Clamp_N20N0D
.SUBCKT sg13g2_Clamp_N20N0D
* device instance $1 r0 *1 25.52,4.95 sg13_hv_nmos
M$1 sub! \$5 \$6 sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $2 r0 *1 27.3,4.95 sg13_hv_nmos
M$2 \$6 \$5 sub! sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $3 r0 *1 28.54,4.95 sg13_hv_nmos
M$3 sub! \$5 \$7 sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $4 r0 *1 30.32,4.95 sg13_hv_nmos
M$4 \$7 \$5 sub! sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $5 r0 *1 31.56,4.95 sg13_hv_nmos
M$5 sub! \$5 \$8 sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $6 r0 *1 33.34,4.95 sg13_hv_nmos
M$6 \$8 \$5 sub! sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $7 r0 *1 34.58,4.95 sg13_hv_nmos
M$7 sub! \$5 \$9 sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $8 r0 *1 36.36,4.95 sg13_hv_nmos
M$8 \$9 \$5 sub! sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $9 r0 *1 37.6,4.95 sg13_hv_nmos
M$9 sub! \$5 \$10 sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $10 r0 *1 39.38,4.95 sg13_hv_nmos
M$10 \$10 \$5 sub! sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $11 r0 *1 40.62,4.95 sg13_hv_nmos
M$11 sub! \$5 \$11 sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $12 r0 *1 42.4,4.95 sg13_hv_nmos
M$12 \$11 \$5 sub! sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $13 r0 *1 43.64,4.95 sg13_hv_nmos
M$13 sub! \$5 \$12 sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $14 r0 *1 45.42,4.95 sg13_hv_nmos
M$14 \$12 \$5 sub! sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $15 r0 *1 46.66,4.95 sg13_hv_nmos
M$15 sub! \$5 \$13 sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $16 r0 *1 48.44,4.95 sg13_hv_nmos
M$16 \$13 \$5 sub! sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $17 r0 *1 49.68,4.95 sg13_hv_nmos
M$17 sub! \$5 \$14 sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $18 r0 *1 51.46,4.95 sg13_hv_nmos
M$18 \$14 \$5 sub! sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $19 r0 *1 52.7,4.95 sg13_hv_nmos
M$19 sub! \$5 \$15 sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $20 r0 *1 54.48,4.95 sg13_hv_nmos
M$20 \$15 \$5 sub! sub! sg13_hv_nmos W=4.3999999999999995 L=0.5999999999999998
* device instance $21 r0 *1 66.305,2.75 rppd
R$21 sub! \$5 rppd w=0.5 l=3.54 ps=0 b=0 m=1
.ENDS sg13g2_Clamp_N20N0D

* Extracted by KLayout with SG13G2 LVS runset on : 10/05/2024 21:06

* cell UHEE628_S2024
* pin PAD,RES
* pin CK4,PAD
* pin CK5,PAD
* pin CK6,PAD
* pin IOVDD
* pin AVDD
* pin CORE
* pin CORE
* pin CORE
* pin CORE
* pin IN6,PAD
* pin OUT6
* pin VDD
* pin dout
* pin CORE
* pin IN5,PAD
* pin OUT5
* pin CORE
* pin IN4,PAD
* pin OUT4
* pin CORE
* pin PAD,VLO
* pin CORE
* pin PAD,VHI
* pin CORE
* pin IN3,PAD
* pin OUT3
* pin CORE
* pin PAD,VLDO
* pin IN2,PAD
* pin OUT2
* pin CORE
* pin CORE
* pin IN1,PAD
* pin OUT1
* pin CORE
* pin PAD,VREF
* pin CORE
* pin CORE
* pin CORE
* pin CORE
* pin CK3,PAD
* pin CK2,PAD
* pin CK1,PAD
* pin VSS
.SUBCKT UHEE628_S2024 PAD|RES CK4|PAD CK5|PAD CK6|PAD IOVDD AVDD CORE CORE$1
+ CORE$2 CORE$3 IN6|PAD OUT6 VDD dout CORE$4 IN5|PAD OUT5 CORE$5 IN4|PAD OUT4
+ CORE$6 PAD|VLO CORE$7 PAD|VHI CORE$8 IN3|PAD OUT3 CORE$9 PAD|VLDO IN2|PAD
+ OUT2 CORE$10 CORE$11 IN1|PAD OUT1 CORE$12 PAD|VREF CORE$13 CORE$14 CORE$15
+ CORE$16 CK3|PAD CK2|PAD CK1|PAD VSS
* device instance $1 r0 *1 500.255,239.005 sg13_lv_nmos
M$1 \$4796 \$4801 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $2 r0 *1 700.255,239.005 sg13_lv_nmos
M$2 \$4797 \$4802 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $3 r0 *1 800.255,239.005 sg13_lv_nmos
M$3 \$4798 \$4803 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $4 r0 *1 900.255,239.005 sg13_lv_nmos
M$4 \$4799 \$4804 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $5 r0 *1 431.875,301.115 sg13_lv_nmos
M$5 \$5939 \$6129 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $7 r0 *1 432.905,301.115 sg13_lv_nmos
M$7 \$5939 \$6407 \$6116 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $9 r0 *1 434.755,301.115 sg13_lv_nmos
M$9 \$5940 \$6130 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $11 r0 *1 435.785,301.115 sg13_lv_nmos
M$11 \$5940 \$6170 \$5941 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $13 r0 *1 437.56,301.14 sg13_lv_nmos
M$13 VSS \$6116 \$5942 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $17 r0 *1 440.44,301.14 sg13_lv_nmos
M$17 VSS \$5941 \$5943 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $21 r0 *1 443.26,301.14 sg13_lv_nmos
M$21 VSS \$5942 \$5944 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $29 r0 *1 448.06,301.14 sg13_lv_nmos
M$29 VSS \$5943 \$5945 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $37 r0 *1 1060.995,297.48 sg13_lv_nmos
M$37 \$5741 dout VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $38 r0 *1 456.79,303.21 sg13_lv_nmos
M$38 VSS \$5945 \$6138 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $39 r0 *1 460.28,303.305 sg13_lv_nmos
M$39 VSS \$5926 \$6143 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $40 r0 *1 461.13,303.21 sg13_lv_nmos
M$40 VSS \$5944 \$6148 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $41 r0 *1 461.44,303.21 sg13_lv_nmos
M$41 \$6148 \$6143 \$6140 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $42 r0 *1 1060.995,300.99 sg13_lv_nmos
M$42 \$5946 dout VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $43 r0 *1 431.085,305.825 sg13_lv_nmos
M$43 VSS \$4799 \$6165 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $45 r0 *1 433.06,305.8 sg13_lv_nmos
M$45 \$6166 \$6165 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $47 r0 *1 434.09,305.8 sg13_lv_nmos
M$47 \$6166 \$6129 \$6178 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $49 r0 *1 435.865,305.825 sg13_lv_nmos
M$49 VSS \$6178 \$6167 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $53 r0 *1 438.745,305.825 sg13_lv_nmos
M$53 VSS \$6167 \$6168 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $57 r0 *1 441.625,305.825 sg13_lv_nmos
M$57 VSS \$6168 \$6169 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $61 r0 *1 444.505,305.825 sg13_lv_nmos
M$61 VSS \$6169 \$6170 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $65 r0 *1 447.385,305.825 sg13_lv_nmos
M$65 VSS \$6170 \$6171 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $69 r0 *1 450.265,305.825 sg13_lv_nmos
M$69 VSS \$6171 \$6130 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $73 r0 *1 457.97,303.37 sg13_lv_nmos
M$73 \$6142 \$5944 \$6157 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $74 r0 *1 458.48,303.37 sg13_lv_nmos
M$74 VSS \$5926 \$6157 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $75 r0 *1 458.99,303.32 sg13_lv_nmos
M$75 VSS \$6142 \$6139 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $76 r0 *1 465.4,304.425 sg13_lv_nmos
M$76 \$6144 \$6171 \$6133 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $77 r0 *1 465.91,304.425 sg13_lv_nmos
M$77 \$6133 \$5944 \$6145 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $78 r0 *1 469.22,304.415 sg13_lv_nmos
M$78 \$6118 \$5945 \$6145 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $79 r0 *1 469.73,304.415 sg13_lv_nmos
M$79 \$6145 \$4796 \$6117 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $80 r0 *1 431.05,310.465 sg13_lv_nmos
M$80 VSS \$6165 \$6402 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $82 r0 *1 433.025,310.44 sg13_lv_nmos
M$82 \$6212 \$6130 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $84 r0 *1 434.055,310.44 sg13_lv_nmos
M$84 \$6212 \$6402 \$6403 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $86 r0 *1 435.83,310.475 sg13_lv_nmos
M$86 VSS \$6403 \$6404 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $90 r0 *1 438.71,310.475 sg13_lv_nmos
M$90 VSS \$6404 \$6405 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $94 r0 *1 441.59,310.475 sg13_lv_nmos
M$94 VSS \$6405 \$6406 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $98 r0 *1 444.47,310.475 sg13_lv_nmos
M$98 VSS \$6406 \$6407 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $102 r0 *1 447.35,310.475 sg13_lv_nmos
M$102 VSS \$6407 \$6408 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $106 r0 *1 450.23,310.475 sg13_lv_nmos
M$106 VSS \$6408 \$6129 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $110 r0 *1 457.825,307.85 sg13_lv_nmos
M$110 \$6193 \$6139 PAD|VLO VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $111 r0 *1 460.21,307.855 sg13_lv_nmos
M$111 \$6193 \$5945 \$6197 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $112 r0 *1 465.395,308.555 sg13_lv_nmos
M$112 VSS \$6144 \$6144 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $113 r0 *1 469.615,308.555 sg13_lv_nmos
M$113 VSS \$6118 \$6117 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $114 r0 *1 431.685,321.635 sg13_lv_nmos
M$114 VSS \$5944 \$6971 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $115 r0 *1 432.865,321.795 sg13_lv_nmos
M$115 \$6972 \$5945 \$7042 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $116 r0 *1 433.375,321.795 sg13_lv_nmos
M$116 VSS \$6782 \$7042 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $117 r0 *1 433.885,321.745 sg13_lv_nmos
M$117 VSS \$6972 \$6973 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $118 r0 *1 435.175,321.73 sg13_lv_nmos
M$118 VSS \$6782 \$6974 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $119 r0 *1 436.025,321.635 sg13_lv_nmos
M$119 VSS \$5945 \$7045 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $120 r0 *1 436.335,321.635 sg13_lv_nmos
M$120 \$7045 \$6974 \$6975 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $121 r0 *1 440.295,322.85 sg13_lv_nmos
M$121 \$7039 \$6408 \$6774 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $122 r0 *1 440.805,322.85 sg13_lv_nmos
M$122 \$6774 \$5945 \$7040 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $123 r0 *1 444.115,322.84 sg13_lv_nmos
M$123 \$6783 \$5944 \$7040 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $124 r0 *1 444.625,322.84 sg13_lv_nmos
M$124 \$7040 \$4796 \$6197 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $125 r0 *1 451.1,325.71 sg13_lv_nmos
M$125 VSS \$5944 \$7301 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $126 r0 *1 452.54,325.71 sg13_lv_nmos
M$126 VSS \$4796 \$7302 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $127 r0 *1 453.94,325.71 sg13_lv_nmos
M$127 VSS \$7322 \$5926 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $129 r0 *1 454.96,325.76 sg13_lv_nmos
M$129 VSS \$7385 \$7322 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $130 r0 *1 456.195,325.53 sg13_lv_nmos
M$130 \$7303 \$7385 \$7321 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $131 r0 *1 456.505,325.53 sg13_lv_nmos
M$131 \$7321 \$7302 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $132 r0 *1 457.085,325.915 sg13_lv_nmos
M$132 VSS \$7323 \$7304 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $133 r0 *1 464.925,325.53 sg13_lv_nmos
M$133 \$7306 \$7307 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $134 r0 *1 465.435,325.53 sg13_lv_nmos
M$134 VSS \$7302 \$7318 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $135 r0 *1 465.745,325.53 sg13_lv_nmos
M$135 \$7318 \$7316 \$7307 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $136 r0 *1 467.785,325.64 sg13_lv_nmos
M$136 VSS \$7316 \$7309 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $137 r0 *1 466.765,325.69 sg13_lv_nmos
M$137 VSS \$7316 \$7308 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $139 r0 *1 468.805,325.69 sg13_lv_nmos
M$139 VSS \$7309 \$6782 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $141 r0 *1 470.56,325.71 sg13_lv_nmos
M$141 VSS \$6782 dout VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $143 r0 *1 432.72,326.275 sg13_lv_nmos
M$143 \$7314 \$6973 PAD|VLO VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $144 r0 *1 435.105,326.28 sg13_lv_nmos
M$144 \$7314 \$5944 CORE$4 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $145 r0 *1 440.29,326.98 sg13_lv_nmos
M$145 VSS \$7039 \$7039 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $146 r0 *1 444.51,326.98 sg13_lv_nmos
M$146 VSS \$6783 \$6197 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $147 r0 *1 457.62,331.325 sg13_lv_nmos
M$147 \$7364 \$5944 \$6117 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $148 r0 *1 458.175,325.595 sg13_lv_nmos
M$148 VSS \$7302 \$7320 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $149 r0 *1 458.485,325.595 sg13_lv_nmos
M$149 \$7320 \$7304 \$7315 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $150 r0 *1 459.26,326.32 sg13_lv_nmos
M$150 \$7303 \$7305 \$7323 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $151 r0 *1 459.77,326.32 sg13_lv_nmos
M$151 \$7323 \$7339 \$7315 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $152 r0 *1 460.575,329.87 sg13_lv_nmos
M$152 VSS \$6144 \$7371 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $153 r0 *1 460.575,330.815 sg13_lv_nmos
M$153 \$7371 \$5945 \$7377 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $154 r0 *1 460.575,331.325 sg13_lv_nmos
M$154 \$7377 \$7378 \$7383 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $155 r0 *1 461.03,325.795 sg13_lv_nmos
M$155 VSS \$7305 \$7339 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $156 r0 *1 462.13,325.795 sg13_lv_nmos
M$156 VSS \$5944 \$7305 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $157 r0 *1 463.65,329.87 sg13_lv_nmos
M$157 VSS \$7364 \$7372 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $158 r0 *1 463.65,330.815 sg13_lv_nmos
M$158 \$7372 \$5945 \$7379 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $159 r0 *1 463.65,331.325 sg13_lv_nmos
M$159 \$7379 \$7383 \$7378 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $160 r0 *1 463.34,325.915 sg13_lv_nmos
M$160 \$7316 \$7305 \$7306 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $161 r0 *1 463.875,325.755 sg13_lv_nmos
M$161 \$7304 \$7339 \$7316 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $162 r0 *1 467.385,330.81 sg13_lv_nmos
M$162 VSS \$7378 \$7380 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $163 r0 *1 467.385,331.32 sg13_lv_nmos
M$163 \$7380 \$7385 \$7384 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $164 r0 *1 470.52,330.81 sg13_lv_nmos
M$164 VSS \$7383 \$7381 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $165 r0 *1 470.52,331.32 sg13_lv_nmos
M$165 \$7381 \$7384 \$7385 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $166 r0 *1 458.328,399.377 sg13_lv_nmos
M$166 \$9634 \$9658 CORE$5 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $167 r0 *1 459.485,394.652 sg13_lv_nmos
M$167 PAD|VLO \$9628 \$9634 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $168 r0 *1 464.231,393.708 sg13_lv_nmos
M$168 \$9628 \$9632 VSS VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $169 r0 *1 464.741,393.758 sg13_lv_nmos
M$169 VSS \$9659 \$9637 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $170 r0 *1 465.251,393.758 sg13_lv_nmos
M$170 \$9637 \$10180 \$9632 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $171 r0 *1 476.371,393.758 sg13_lv_nmos
M$171 \$9633 \$9658 \$9639 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $172 r0 *1 476.881,393.758 sg13_lv_nmos
M$172 VSS \$9635 \$9639 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $173 r0 *1 477.391,393.708 sg13_lv_nmos
M$173 VSS \$9633 \$9629 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $174 r0 *1 482.137,394.652 sg13_lv_nmos
M$174 PAD|VLO \$9629 \$9848 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $175 r0 *1 483.294,399.377 sg13_lv_nmos
M$175 \$10410 \$10180 \$9848 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $176 r0 *1 1060.995,397.48 sg13_lv_nmos
M$176 \$9650 \$9659 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $177 r0 *1 1060.995,400.99 sg13_lv_nmos
M$177 \$10174 \$9659 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $178 r0 *1 443.526,403.27 sg13_lv_nmos
M$178 \$10369 \$10180 \$9623 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $179 r0 *1 448.102,403.27 sg13_lv_nmos
M$179 \$9623 \$11334 \$10183 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $180 r0 *1 493.52,403.27 sg13_lv_nmos
M$180 \$10184 \$10931 \$9624 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $181 r0 *1 498.096,403.27 sg13_lv_nmos
M$181 \$9624 \$9658 \$10370 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $182 r0 *1 454.041,411.248 sg13_lv_nmos
M$182 \$10183 \$10183 VSS VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $183 r0 *1 458.723,405.86 sg13_lv_nmos
M$183 VSS \$9658 \$9842 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $184 r0 *1 462.071,405.955 sg13_lv_nmos
M$184 VSS \$9659 \$10208 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $185 r0 *1 462.921,405.86 sg13_lv_nmos
M$185 VSS \$10180 \$10214 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $186 r0 *1 463.231,405.86 sg13_lv_nmos
M$186 \$10214 \$10208 \$10206 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $187 r0 *1 478.391,405.86 sg13_lv_nmos
M$187 \$10207 \$10209 \$10216 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $188 r0 *1 478.701,405.86 sg13_lv_nmos
M$188 \$10216 \$9658 VSS VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $189 r0 *1 479.551,405.955 sg13_lv_nmos
M$189 VSS \$9635 \$10209 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $190 r0 *1 482.899,405.86 sg13_lv_nmos
M$190 \$9843 \$10180 VSS VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $191 r0 *1 487.581,411.248 sg13_lv_nmos
M$191 VSS \$10184 \$10184 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $192 r0 *1 454.041,420.794 sg13_lv_nmos
M$192 \$10410 \$9622 VSS VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $193 r0 *1 458.979,423.251 sg13_lv_nmos
M$193 \$10410 \$4796 \$10369 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $194 r0 *1 463.555,423.251 sg13_lv_nmos
M$194 \$10369 \$9658 \$9622 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $195 r0 *1 478.067,423.251 sg13_lv_nmos
M$195 \$9625 \$10180 \$10370 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $196 r0 *1 482.643,423.251 sg13_lv_nmos
M$196 \$10370 \$4796 \$10411 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $197 r0 *1 487.581,420.794 sg13_lv_nmos
M$197 VSS \$9625 \$10411 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $198 r0 *1 452.732,430.97 sg13_lv_nmos
M$198 \$10925 \$11326 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $200 r0 *1 453.762,430.97 sg13_lv_nmos
M$200 \$10925 \$11335 \$10926 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $202 r0 *1 455.996,430.995 sg13_lv_nmos
M$202 VSS \$10926 \$10927 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $206 r0 *1 459.411,430.995 sg13_lv_nmos
M$206 VSS \$10927 \$10928 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $210 r0 *1 462.647,430.995 sg13_lv_nmos
M$210 VSS \$10928 \$10929 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $214 r0 *1 466.172,430.995 sg13_lv_nmos
M$214 VSS \$10929 \$10930 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $218 r0 *1 470.029,430.995 sg13_lv_nmos
M$218 VSS \$10930 \$10931 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $222 r0 *1 473.998,430.995 sg13_lv_nmos
M$222 VSS \$10931 \$10932 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $226 r0 *1 477.918,430.97 sg13_lv_nmos
M$226 \$10933 \$10932 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $228 r0 *1 478.948,430.97 sg13_lv_nmos
M$228 \$10933 \$10930 \$10934 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $230 r0 *1 481.602,430.995 sg13_lv_nmos
M$230 VSS \$10934 \$10935 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $234 r0 *1 484.998,430.995 sg13_lv_nmos
M$234 VSS \$10935 \$10180 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $242 r0 *1 446.843,438.963 sg13_lv_nmos
M$242 VSS \$4798 \$11326 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $244 r0 *1 449.364,438.963 sg13_lv_nmos
M$244 VSS \$11326 \$11327 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $246 r0 *1 452.01,438.938 sg13_lv_nmos
M$246 \$11328 \$11327 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $248 r0 *1 453.04,438.938 sg13_lv_nmos
M$248 \$11328 \$10932 \$11329 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $250 r0 *1 455.373,438.964 sg13_lv_nmos
M$250 VSS \$11329 \$11330 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $254 r0 *1 459.841,438.964 sg13_lv_nmos
M$254 VSS \$11330 \$11331 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $258 r0 *1 463.257,438.964 sg13_lv_nmos
M$258 VSS \$11331 \$11332 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $262 r0 *1 466.777,438.964 sg13_lv_nmos
M$262 VSS \$11332 \$11333 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $266 r0 *1 470.634,438.964 sg13_lv_nmos
M$266 VSS \$11333 \$11334 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $270 r0 *1 474.603,438.964 sg13_lv_nmos
M$270 VSS \$11334 \$11335 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $274 r0 *1 478.273,438.939 sg13_lv_nmos
M$274 \$11336 \$11335 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $276 r0 *1 479.303,438.939 sg13_lv_nmos
M$276 \$11336 \$11333 \$11337 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $278 r0 *1 480.059,445.671 sg13_lv_nmos
M$278 VSS \$11659 \$11517 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $279 r0 *1 481.957,438.964 sg13_lv_nmos
M$279 VSS \$11337 \$11338 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $283 r0 *1 485.353,438.964 sg13_lv_nmos
M$283 VSS \$11338 \$9658 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $291 r0 *1 450.192,450.371 sg13_lv_nmos
M$291 VSS \$11690 \$11713 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $292 r0 *1 449.324,446.442 sg13_lv_nmos
M$292 VSS \$11666 \$9635 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $294 r0 *1 450.344,446.492 sg13_lv_nmos
M$294 VSS \$11717 \$11666 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $295 r0 *1 452.324,446.262 sg13_lv_nmos
M$295 \$11649 \$11717 \$11672 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $296 r0 *1 452.634,446.262 sg13_lv_nmos
M$296 \$11672 \$11650 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $297 r0 *1 453.214,446.647 sg13_lv_nmos
M$297 VSS \$11686 \$11651 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $298 r0 *1 454.304,446.327 sg13_lv_nmos
M$298 VSS \$11650 \$11673 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $299 r0 *1 454.614,446.327 sg13_lv_nmos
M$299 \$11673 \$11651 \$11652 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $300 r0 *1 455.389,447.052 sg13_lv_nmos
M$300 \$11649 \$11653 \$11686 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $301 r0 *1 455.899,447.052 sg13_lv_nmos
M$301 \$11686 \$11667 \$11652 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $302 r0 *1 457.159,446.527 sg13_lv_nmos
M$302 VSS \$11653 \$11667 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $303 r0 *1 458.259,446.527 sg13_lv_nmos
M$303 VSS \$9658 \$11653 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $304 r0 *1 459.469,446.647 sg13_lv_nmos
M$304 \$11668 \$11653 \$11654 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $305 r0 *1 460.004,446.487 sg13_lv_nmos
M$305 \$11651 \$11667 \$11668 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $306 r0 *1 461.054,446.262 sg13_lv_nmos
M$306 \$11654 \$11655 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $307 r0 *1 461.564,446.262 sg13_lv_nmos
M$307 VSS \$11650 \$11677 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $308 r0 *1 461.874,446.262 sg13_lv_nmos
M$308 \$11677 \$11668 \$11655 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $309 r0 *1 463.914,446.372 sg13_lv_nmos
M$309 VSS \$11668 \$11657 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $310 r0 *1 462.894,446.422 sg13_lv_nmos
M$310 VSS \$11668 \$11656 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $312 r0 *1 464.934,446.422 sg13_lv_nmos
M$312 VSS \$11657 \$9659 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $314 r0 *1 467.705,446.442 sg13_lv_nmos
M$314 VSS \$4796 \$11650 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $315 r0 *1 469.14,446.442 sg13_lv_nmos
M$315 VSS \$9658 \$11658 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $316 r0 *1 469.693,451.053 sg13_lv_nmos
M$316 \$11659 \$9658 \$10411 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $317 r0 *1 480.059,451.332 sg13_lv_nmos
M$317 VSS \$10184 \$11706 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $318 r0 *1 483.419,452.999 sg13_lv_nmos
M$318 \$11690 \$11646 \$11718 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $319 r0 *1 483.419,447.338 sg13_lv_nmos
M$319 \$11646 \$11690 \$11669 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $320 r0 *1 485.064,447.338 sg13_lv_nmos
M$320 \$11669 \$10180 \$11517 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $321 r0 *1 485.064,452.999 sg13_lv_nmos
M$321 \$11718 \$10180 \$11706 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $322 r0 *1 450.192,456.171 sg13_lv_nmos
M$322 VSS \$11646 \$12328 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $323 r0 *1 450.234,459.67 sg13_lv_nmos
M$323 \$12329 \$11717 \$12328 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $324 r0 *1 450.234,453.87 sg13_lv_nmos
M$324 \$11717 \$12329 \$11713 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $325 r0 *1 1060.995,497.48 sg13_lv_nmos
M$325 \$13602 \$13736 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $326 r0 *1 1060.995,500.99 sg13_lv_nmos
M$326 \$13982 \$13736 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $327 r0 *1 485.618,504.427 sg13_lv_nmos
M$327 \$14006 \$14016 \$14026 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $328 r0 *1 486.008,504.427 sg13_lv_nmos
M$328 \$14026 \$14007 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $329 r0 *1 486.568,504.427 sg13_lv_nmos
M$329 VSS \$13993 \$14020 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $330 r0 *1 486.923,504.427 sg13_lv_nmos
M$330 \$14020 \$14006 \$14007 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $331 r0 *1 483.978,504.537 sg13_lv_nmos
M$331 VSS \$14004 \$14005 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $332 r0 *1 484.648,504.537 sg13_lv_nmos
M$332 \$14005 \$13999 \$14006 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $333 r0 *1 482.098,504.652 sg13_lv_nmos
M$333 \$14003 \$14016 \$14004 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $334 r0 *1 482.608,504.652 sg13_lv_nmos
M$334 \$14004 \$13999 \$14025 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $335 r0 *1 482.998,504.652 sg13_lv_nmos
M$335 \$14025 \$14005 \$14024 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $336 r0 *1 483.358,504.652 sg13_lv_nmos
M$336 VSS \$13993 \$14024 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $337 r0 *1 476.768,504.592 sg13_lv_nmos
M$337 VSS \$14713 \$14002 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $338 r0 *1 478.818,504.452 sg13_lv_nmos
M$338 \$14003 \$14233 \$14029 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $339 r0 *1 479.188,504.452 sg13_lv_nmos
M$339 \$14029 \$13993 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $340 r0 *1 487.963,504.592 sg13_lv_nmos
M$340 VSS \$14006 \$14008 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $341 r0 *1 489.163,504.497 sg13_lv_nmos
M$341 \$14009 \$14006 VSS VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $342 r0 *1 489.703,504.592 sg13_lv_nmos
M$342 VSS \$14009 \$14010 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $343 r0 *1 491.898,504.592 sg13_lv_nmos
M$343 VSS \$14010 \$13736 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $345 r0 *1 494.693,504.591 sg13_lv_nmos
M$345 VSS \$4796 \$13993 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $346 r0 *1 496.608,504.591 sg13_lv_nmos
M$346 VSS \$14030 \$14011 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $348 r0 *1 497.628,504.641 sg13_lv_nmos
M$348 VSS \$14233 \$14030 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $349 r0 *1 480.333,504.767 sg13_lv_nmos
M$349 VSS \$14713 \$14016 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $350 r0 *1 480.843,504.767 sg13_lv_nmos
M$350 VSS \$14016 \$13999 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $351 r0 *1 481.503,510.997 sg13_lv_nmos
M$351 VSS \$14194 \$14199 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $352 r0 *1 483.503,509.467 sg13_lv_nmos
M$352 \$14121 \$14713 \$14122 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $353 r0 *1 485.503,510.997 sg13_lv_nmos
M$353 VSS \$14122 \$14200 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $354 r0 *1 438.155,518.846 sg13_lv_nmos
M$354 VSS \$14241 \$14242 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $358 r0 *1 441.035,518.846 sg13_lv_nmos
M$358 VSS \$14242 \$14243 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $362 r0 *1 443.915,518.846 sg13_lv_nmos
M$362 VSS \$14243 \$14244 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $366 r0 *1 446.795,518.846 sg13_lv_nmos
M$366 VSS \$14244 \$14245 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $370 r0 *1 449.675,518.846 sg13_lv_nmos
M$370 VSS \$14245 \$14246 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $374 r0 *1 452.555,518.846 sg13_lv_nmos
M$374 VSS \$14246 \$14247 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $378 r0 *1 458.315,518.846 sg13_lv_nmos
M$378 VSS \$14248 \$14249 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $382 r0 *1 461.135,518.846 sg13_lv_nmos
M$382 VSS \$14249 \$14250 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $390 r0 *1 481.703,513.099 sg13_lv_nmos
M$390 \$14199 \$14250 \$14205 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $391 r0 *1 482.903,513.099 sg13_lv_nmos
M$391 \$14205 \$14232 \$14206 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $392 r0 *1 484.103,513.099 sg13_lv_nmos
M$392 \$14232 \$14206 \$14207 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $393 r0 *1 485.303,513.099 sg13_lv_nmos
M$393 \$14207 \$14250 \$14200 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $394 r0 *1 488.561,513.099 sg13_lv_nmos
M$394 VSS \$14232 \$14208 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $395 r0 *1 489.761,513.099 sg13_lv_nmos
M$395 \$14208 \$14233 \$14209 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $396 r0 *1 490.961,513.099 sg13_lv_nmos
M$396 \$14233 \$14209 \$14210 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $397 r0 *1 492.161,513.099 sg13_lv_nmos
M$397 \$14210 \$14206 VSS VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $398 r0 *1 431.455,521.281 sg13_lv_nmos
M$398 VSS \$4797 \$14258 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $400 r0 *1 433.375,521.281 sg13_lv_nmos
M$400 VSS \$14258 \$14702 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $402 r0 *1 435.35,518.871 sg13_lv_nmos
M$402 \$14271 \$14709 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $404 r0 *1 436.38,518.871 sg13_lv_nmos
M$404 \$14271 \$14258 \$14241 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $406 r0 *1 435.35,521.256 sg13_lv_nmos
M$406 \$14703 \$14247 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $408 r0 *1 436.38,521.256 sg13_lv_nmos
M$408 \$14703 \$14702 \$14718 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $410 r0 *1 438.155,521.281 sg13_lv_nmos
M$410 VSS \$14718 \$14704 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $414 r0 *1 441.035,521.281 sg13_lv_nmos
M$414 VSS \$14704 \$14705 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $418 r0 *1 443.915,521.281 sg13_lv_nmos
M$418 VSS \$14705 \$14706 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $422 r0 *1 446.795,521.281 sg13_lv_nmos
M$422 VSS \$14706 \$14707 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $426 r0 *1 449.675,521.281 sg13_lv_nmos
M$426 VSS \$14707 \$14708 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $430 r0 *1 452.555,521.281 sg13_lv_nmos
M$430 VSS \$14708 \$14709 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $434 r0 *1 455.51,518.871 sg13_lv_nmos
M$434 \$14272 \$14247 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $436 r0 *1 456.54,518.871 sg13_lv_nmos
M$436 \$14272 \$14245 \$14248 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $438 r0 *1 455.51,521.256 sg13_lv_nmos
M$438 \$14710 \$14709 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $440 r0 *1 456.54,521.256 sg13_lv_nmos
M$440 \$14710 \$14707 \$14711 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $442 r0 *1 458.315,521.281 sg13_lv_nmos
M$442 VSS \$14711 \$14712 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $446 r0 *1 461.135,521.281 sg13_lv_nmos
M$446 VSS \$14712 \$14713 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $454 r0 *1 431.5,535.261 sg13_lv_nmos
M$454 VSS \$14713 \$15026 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $455 r0 *1 432.935,535.356 sg13_lv_nmos
M$455 VSS \$14010 \$15033 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $456 r0 *1 433.785,535.261 sg13_lv_nmos
M$456 VSS \$14250 \$15038 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $457 r0 *1 434.095,535.261 sg13_lv_nmos
M$457 \$15038 \$15033 \$15027 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $458 r0 *1 435.785,535.421 sg13_lv_nmos
M$458 \$15034 \$14250 \$15040 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $459 r0 *1 436.295,535.421 sg13_lv_nmos
M$459 VSS \$14010 \$15040 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $460 r0 *1 436.805,535.371 sg13_lv_nmos
M$460 VSS \$15034 \$15028 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $461 r0 *1 443.55,535.276 sg13_lv_nmos
M$461 VSS \$15029 \$15029 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $462 r0 *1 455.2,535.261 sg13_lv_nmos
M$462 VSS \$15047 \$15048 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $463 r0 *1 466.5,535.261 sg13_lv_nmos
M$463 VSS \$14250 \$15030 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $464 r0 *1 467.935,535.356 sg13_lv_nmos
M$464 VSS \$14011 \$15035 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $465 r0 *1 468.785,535.261 sg13_lv_nmos
M$465 VSS \$14713 \$15044 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $466 r0 *1 469.095,535.261 sg13_lv_nmos
M$466 \$15044 \$15035 \$15031 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $467 r0 *1 470.785,535.421 sg13_lv_nmos
M$467 \$15036 \$14713 \$15046 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $468 r0 *1 471.295,535.421 sg13_lv_nmos
M$468 VSS \$14011 \$15046 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $469 r0 *1 471.805,535.371 sg13_lv_nmos
M$469 VSS \$15036 \$15032 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $470 r0 *1 478.55,535.276 sg13_lv_nmos
M$470 VSS \$14194 \$14194 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $471 r0 *1 490.2,535.261 sg13_lv_nmos
M$471 VSS \$15049 \$14121 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $472 r0 *1 454.14,553.166 sg13_lv_nmos
M$472 \$15333 \$14250 \$15341 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $473 r0 *1 455.45,553.166 sg13_lv_nmos
M$473 \$15341 \$14713 \$15047 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $474 r0 *1 456.763,553.166 sg13_lv_nmos
M$474 \$15341 \$4796 \$15048 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $475 r0 *1 489.14,553.166 sg13_lv_nmos
M$475 \$15334 \$14713 \$15335 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $476 r0 *1 490.45,553.166 sg13_lv_nmos
M$476 \$15335 \$14250 \$15049 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $477 r0 *1 491.763,553.166 sg13_lv_nmos
M$477 \$15335 \$4796 \$14121 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $478 r0 *1 434.07,553.206 sg13_lv_nmos
M$478 \$15336 \$15028 PAD|VLO VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $479 r0 *1 436.815,553.216 sg13_lv_nmos
M$479 \$15336 \$14713 CORE$6 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $480 r0 *1 444.09,553.171 sg13_lv_nmos
M$480 \$15029 \$14708 \$15333 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $481 r0 *1 469.07,553.206 sg13_lv_nmos
M$481 \$15076 \$15032 PAD|VLO VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $482 r0 *1 471.815,553.216 sg13_lv_nmos
M$482 \$15076 \$14250 \$15048 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $483 r0 *1 479.09,553.171 sg13_lv_nmos
M$483 \$14194 \$14246 \$15334 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $484 r0 *1 449.83,597.155 sg13_lv_nmos
M$484 \$16921 \$17062 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $486 r0 *1 450.86,597.155 sg13_lv_nmos
M$486 \$16921 \$16931 \$16932 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $488 r0 *1 469.99,597.155 sg13_lv_nmos
M$488 \$16928 \$16927 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $490 r0 *1 471.02,597.155 sg13_lv_nmos
M$490 \$16928 \$16925 \$16933 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $492 r0 *1 452.635,597.18 sg13_lv_nmos
M$492 VSS \$16932 \$16922 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $496 r0 *1 455.515,597.18 sg13_lv_nmos
M$496 VSS \$16922 \$16923 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $500 r0 *1 458.395,597.18 sg13_lv_nmos
M$500 VSS \$16923 \$16924 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $504 r0 *1 461.275,597.18 sg13_lv_nmos
M$504 VSS \$16924 \$16925 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $508 r0 *1 464.155,597.18 sg13_lv_nmos
M$508 VSS \$16925 \$16926 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $512 r0 *1 467.035,597.18 sg13_lv_nmos
M$512 VSS \$16926 \$16927 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $516 r0 *1 472.795,597.18 sg13_lv_nmos
M$516 VSS \$16933 \$16929 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $520 r0 *1 475.615,597.18 sg13_lv_nmos
M$520 VSS \$16929 \$16930 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $528 r0 *1 445.935,602.98 sg13_lv_nmos
M$528 VSS \$16829 \$16931 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $530 r0 *1 447.855,602.98 sg13_lv_nmos
M$530 VSS \$16931 \$17055 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $532 r0 *1 449.83,602.955 sg13_lv_nmos
M$532 \$17056 \$16927 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $534 r0 *1 450.86,602.955 sg13_lv_nmos
M$534 \$17056 \$17055 \$17066 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $536 r0 *1 452.635,602.98 sg13_lv_nmos
M$536 VSS \$17066 \$17057 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $540 r0 *1 455.515,602.98 sg13_lv_nmos
M$540 VSS \$17057 \$17058 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $544 r0 *1 458.395,602.98 sg13_lv_nmos
M$544 VSS \$17058 \$17059 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $548 r0 *1 461.275,602.98 sg13_lv_nmos
M$548 VSS \$17059 \$17060 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $552 r0 *1 464.155,602.98 sg13_lv_nmos
M$552 VSS \$17060 \$17061 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $556 r0 *1 467.035,602.98 sg13_lv_nmos
M$556 VSS \$17061 \$17062 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $560 r0 *1 469.99,602.955 sg13_lv_nmos
M$560 \$17063 \$17062 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $562 r0 *1 471.02,602.955 sg13_lv_nmos
M$562 \$17063 \$17060 \$17067 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $564 r0 *1 472.795,602.98 sg13_lv_nmos
M$564 VSS \$17067 \$17064 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $568 r0 *1 475.615,602.98 sg13_lv_nmos
M$568 VSS \$17064 \$17065 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $576 r0 *1 433.27,616.415 sg13_lv_nmos
M$576 VSS \$17065 \$17383 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $577 r0 *1 434.36,616.51 sg13_lv_nmos
M$577 VSS \$17226 \$17384 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $578 r0 *1 435.21,616.415 sg13_lv_nmos
M$578 VSS \$16930 \$17397 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $579 r0 *1 435.52,616.415 sg13_lv_nmos
M$579 \$17397 \$17384 \$17381 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $580 r0 *1 436.85,616.575 sg13_lv_nmos
M$580 \$17388 \$16930 \$17398 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $581 r0 *1 437.36,616.575 sg13_lv_nmos
M$581 VSS \$17226 \$17398 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $582 r0 *1 437.87,616.525 sg13_lv_nmos
M$582 VSS \$17388 \$17369 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $583 r0 *1 441.655,618.475 sg13_lv_nmos
M$583 PAD|VLO \$17369 \$17495 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $584 r0 *1 454.37,616.04 sg13_lv_nmos
M$584 \$17370 \$17061 \$17393 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $585 r0 *1 454.37,616.55 sg13_lv_nmos
M$585 \$17393 \$16930 \$17673 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $586 r0 *1 454.37,617.83 sg13_lv_nmos
M$586 \$17412 \$17065 \$17673 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $587 r0 *1 454.37,618.34 sg13_lv_nmos
M$587 \$17673 \$4796 \$17496 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $588 r0 *1 469.325,616.415 sg13_lv_nmos
M$588 VSS \$16930 \$17385 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $589 r0 *1 470.415,616.51 sg13_lv_nmos
M$589 VSS \$17355 \$17386 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $590 r0 *1 471.265,616.415 sg13_lv_nmos
M$590 VSS \$17065 \$17406 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $591 r0 *1 471.575,616.415 sg13_lv_nmos
M$591 \$17406 \$17386 \$17382 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $592 r0 *1 472.905,616.575 sg13_lv_nmos
M$592 \$17389 \$17065 \$17404 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $593 r0 *1 473.415,616.575 sg13_lv_nmos
M$593 VSS \$17355 \$17404 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $594 r0 *1 473.925,616.525 sg13_lv_nmos
M$594 VSS \$17389 \$17371 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $595 r0 *1 477.71,618.475 sg13_lv_nmos
M$595 PAD|VLO \$17371 \$17540 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $596 r0 *1 490.425,616.04 sg13_lv_nmos
M$596 \$17372 \$16926 \$17394 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $597 r0 *1 490.425,616.55 sg13_lv_nmos
M$597 \$17394 \$17065 \$17674 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $598 r0 *1 490.425,617.83 sg13_lv_nmos
M$598 \$17413 \$16930 \$17674 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $599 r0 *1 490.425,618.34 sg13_lv_nmos
M$599 \$17674 \$4796 \$17497 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $600 r0 *1 505.425,616.53 sg13_lv_nmos
M$600 VSS \$17065 \$17387 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $601 r0 *1 520.915,619.83 sg13_lv_nmos
M$601 \$17541 \$17650 \$17647 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $602 r0 *1 521.225,619.83 sg13_lv_nmos
M$602 \$17647 \$17536 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $603 r0 *1 521.805,620.215 sg13_lv_nmos
M$603 VSS \$17663 \$17542 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $604 r0 *1 522.895,619.895 sg13_lv_nmos
M$604 VSS \$17536 \$17655 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $605 r0 *1 523.205,619.895 sg13_lv_nmos
M$605 \$17655 \$17542 \$17646 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $606 r0 *1 525.75,620.095 sg13_lv_nmos
M$606 VSS \$17543 \$17651 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $607 r0 *1 526.85,620.095 sg13_lv_nmos
M$607 VSS \$17065 \$17543 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $608 r0 *1 528.06,620.215 sg13_lv_nmos
M$608 \$17652 \$17543 \$17544 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $609 r0 *1 528.595,620.055 sg13_lv_nmos
M$609 \$17542 \$17651 \$17652 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $610 r0 *1 529.645,619.83 sg13_lv_nmos
M$610 \$17544 \$17545 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $611 r0 *1 530.155,619.83 sg13_lv_nmos
M$611 VSS \$17536 \$17649 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $612 r0 *1 530.465,619.83 sg13_lv_nmos
M$612 \$17649 \$17652 \$17545 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $613 r0 *1 532.505,619.94 sg13_lv_nmos
M$613 VSS \$17652 \$17547 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $614 r0 *1 531.485,619.99 sg13_lv_nmos
M$614 VSS \$17652 \$17546 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $616 r0 *1 533.525,619.99 sg13_lv_nmos
M$616 VSS \$17547 \$17226 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $618 r0 *1 535.21,620.01 sg13_lv_nmos
M$618 VSS \$17226 \$17418 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $620 r0 *1 537,620.005 sg13_lv_nmos
M$620 \$17536 \$4796 VSS VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $621 r0 *1 433.495,621.675 sg13_lv_nmos
M$621 CORE$9 \$17065 \$17495 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $622 r0 *1 469.55,621.675 sg13_lv_nmos
M$622 \$17496 \$16930 \$17540 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $623 r0 *1 523.98,620.62 sg13_lv_nmos
M$623 \$17541 \$17543 \$17663 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $624 r0 *1 524.49,620.62 sg13_lv_nmos
M$624 \$17663 \$17651 \$17646 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $625 r0 *1 456.64,623.065 sg13_lv_nmos
M$625 VSS \$17412 \$17496 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $626 r0 *1 462.64,623.065 sg13_lv_nmos
M$626 VSS \$17370 \$17370 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $627 r0 *1 492.695,623.065 sg13_lv_nmos
M$627 VSS \$17413 \$17497 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $628 r0 *1 498.695,623.065 sg13_lv_nmos
M$628 VSS \$17372 \$17372 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $629 r0 *1 505.05,623.5 sg13_lv_nmos
M$629 \$17662 \$17065 \$17497 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $630 r0 *1 509.855,627.99 sg13_lv_nmos
M$630 \$17711 \$16930 \$17721 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $631 r0 *1 509.96,626.51 sg13_lv_nmos
M$631 VSS \$17372 \$17711 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $632 r0 *1 514.795,627.99 sg13_lv_nmos
M$632 \$17712 \$16930 \$17722 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $633 r0 *1 514.885,626.51 sg13_lv_nmos
M$633 VSS \$17662 \$17712 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $634 r0 *1 522.75,627.29 sg13_lv_nmos
M$634 VSS \$17900 \$17713 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $635 r0 *1 523.03,628.795 sg13_lv_nmos
M$635 \$17713 \$17650 \$17727 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $636 r0 *1 529.34,628.76 sg13_lv_nmos
M$636 \$17714 \$17727 \$17650 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $637 r0 *1 529.69,627.28 sg13_lv_nmos
M$637 VSS \$17899 \$17714 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $638 r0 *1 532.795,625.47 sg13_lv_nmos
M$638 VSS \$17703 \$17355 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $640 r0 *1 532.845,626.49 sg13_lv_nmos
M$640 VSS \$17650 \$17703 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $641 r0 *1 509.835,629.77 sg13_lv_nmos
M$641 \$17721 \$17900 \$17899 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $642 r0 *1 514.62,629.77 sg13_lv_nmos
M$642 \$17722 \$17899 \$17900 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $643 r0 *1 1060.995,800.99 sg13_lv_nmos
M$643 \$24446 \$17418 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $644 r0 *1 1060.995,797.48 sg13_lv_nmos
M$644 \$24419 \$17418 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $645 r0 *1 633.21,835.705 sg13_lv_nmos
M$645 VSS \$25483 \$25483 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $647 r0 *1 585.345,846.95 sg13_lv_nmos
M$647 \$25848 \$25867 CORE$11 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $649 r0 *1 592.87,846.075 sg13_lv_nmos
M$649 VSS \$25489 \$25833 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $651 r0 *1 606.935,846.95 sg13_lv_nmos
M$651 \$25849 \$26427 \$25833 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $653 r0 *1 614.46,846.075 sg13_lv_nmos
M$653 VSS \$25490 \$25822 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $655 r0 *1 622.76,843.455 sg13_lv_nmos
M$655 VSS \$25483 \$25825 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $657 r0 *1 623.505,845.055 sg13_lv_nmos
M$657 \$25825 \$26427 \$25834 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $659 r0 *1 623.505,846.655 sg13_lv_nmos
M$659 \$25834 \$25838 \$25839 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $661 r0 *1 626.34,843.455 sg13_lv_nmos
M$661 VSS \$25487 \$25826 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $663 r0 *1 626.465,845.055 sg13_lv_nmos
M$663 \$25826 \$26427 \$25835 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $665 r0 *1 626.465,846.655 sg13_lv_nmos
M$665 \$25835 \$25839 \$25838 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $667 r0 *1 630.06,842.755 sg13_lv_nmos
M$667 \$25822 \$25867 \$25487 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $669 r0 *1 632.73,846.655 sg13_lv_nmos
M$669 \$25836 \$25840 \$25850 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $671 r0 *1 632.73,845.055 sg13_lv_nmos
M$671 VSS \$25838 \$25836 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $673 r0 *1 635.69,845.055 sg13_lv_nmos
M$673 VSS \$25839 \$25837 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $675 r0 *1 635.69,846.655 sg13_lv_nmos
M$675 \$25837 \$25850 \$25840 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $677 r0 *1 586.14,851.955 sg13_lv_nmos
M$677 PAD|VLO \$26460 \$25848 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $678 r0 *1 588.475,852.473 sg13_lv_nmos
M$678 \$25485 \$25867 \$25489 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $679 r0 *1 588.475,849.383 sg13_lv_nmos
M$679 \$25485 \$26427 \$25851 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $680 r0 *1 589.55,849.383 sg13_lv_nmos
M$680 \$25851 \$26999 \$25483 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $681 r0 *1 607.73,851.955 sg13_lv_nmos
M$681 PAD|VLO \$26461 \$25849 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $682 r0 *1 610.065,849.383 sg13_lv_nmos
M$682 \$25486 \$25867 \$25852 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $683 r0 *1 610.065,852.473 sg13_lv_nmos
M$683 \$25486 \$26427 \$25490 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $684 r0 *1 611.14,849.383 sg13_lv_nmos
M$684 \$25852 \$26142 \$25483 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $685 r0 *1 620.94,852.345 sg13_lv_nmos
M$685 VSS \$25867 \$25853 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $686 r0 *1 622.38,852.345 sg13_lv_nmos
M$686 VSS \$4796 \$26446 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $687 r0 *1 623.635,852.165 sg13_lv_nmos
M$687 \$26447 \$25840 \$26464 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $688 r0 *1 623.945,852.165 sg13_lv_nmos
M$688 \$26464 \$26446 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $689 r0 *1 624.525,852.55 sg13_lv_nmos
M$689 VSS \$26494 \$26448 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $690 r0 *1 625.615,852.23 sg13_lv_nmos
M$690 VSS \$26446 \$26485 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $691 r0 *1 625.925,852.23 sg13_lv_nmos
M$691 \$26485 \$26448 \$26449 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $692 r0 *1 628.47,852.43 sg13_lv_nmos
M$692 VSS \$26450 \$26497 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $693 r0 *1 629.57,852.43 sg13_lv_nmos
M$693 VSS \$25867 \$26450 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $694 r0 *1 630.78,852.55 sg13_lv_nmos
M$694 \$26480 \$26450 \$26451 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $695 r0 *1 631.315,852.39 sg13_lv_nmos
M$695 \$26448 \$26497 \$26480 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $696 r0 *1 632.365,852.165 sg13_lv_nmos
M$696 \$26451 \$26452 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $697 r0 *1 632.875,852.165 sg13_lv_nmos
M$697 VSS \$26446 \$26463 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $698 r0 *1 633.185,852.165 sg13_lv_nmos
M$698 \$26463 \$26480 \$26452 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $699 r0 *1 635.225,852.275 sg13_lv_nmos
M$699 VSS \$26480 \$26454 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $700 r0 *1 634.205,852.325 sg13_lv_nmos
M$700 VSS \$26480 \$26453 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $702 r0 *1 636.245,852.325 sg13_lv_nmos
M$702 VSS \$26454 \$26920 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $704 r0 *1 637.86,852.395 sg13_lv_nmos
M$704 VSS \$25840 \$26455 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $705 r0 *1 638.37,852.345 sg13_lv_nmos
M$705 VSS \$26455 \$26921 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $707 r0 *1 640.4,852.345 sg13_lv_nmos
M$707 VSS \$26920 \$28308 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $709 r0 *1 594.145,854.805 sg13_lv_nmos
M$709 \$25485 \$4796 \$25833 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $713 r0 *1 615.735,854.805 sg13_lv_nmos
M$713 \$25486 \$4796 \$25822 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $717 r0 *1 617.465,863.425 sg13_lv_nmos
M$717 \$26922 \$26953 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $719 r0 *1 618.495,863.425 sg13_lv_nmos
M$719 \$26922 \$26954 \$26937 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $721 r0 *1 623.374,863.452 sg13_lv_nmos
M$721 VSS \$26923 \$26924 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $725 r0 *1 626.254,863.452 sg13_lv_nmos
M$725 VSS \$26924 \$26925 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $729 r0 *1 626.7,852.955 sg13_lv_nmos
M$729 \$26447 \$26450 \$26494 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $730 r0 *1 627.21,852.955 sg13_lv_nmos
M$730 \$26494 \$26497 \$26449 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $731 r0 *1 629.134,863.452 sg13_lv_nmos
M$731 VSS \$26925 \$26926 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $735 r0 *1 632.714,863.452 sg13_lv_nmos
M$735 VSS \$26926 \$26142 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $739 r0 *1 636.294,863.452 sg13_lv_nmos
M$739 VSS \$26142 \$26927 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $743 r0 *1 640.7,863.425 sg13_lv_nmos
M$743 \$26928 \$26927 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $745 r0 *1 641.73,863.425 sg13_lv_nmos
M$745 \$26928 \$26926 \$26938 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $747 r0 *1 643.75,863.45 sg13_lv_nmos
M$747 VSS \$26938 \$26929 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $751 r0 *1 646.57,863.452 sg13_lv_nmos
M$751 VSS \$26929 \$26427 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $759 r0 *1 577.495,864.355 sg13_lv_nmos
M$759 \$26956 \$26427 \$26966 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $760 r0 *1 578.005,864.355 sg13_lv_nmos
M$760 VSS \$26920 \$26966 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $761 r0 *1 578.515,864.305 sg13_lv_nmos
M$761 VSS \$26956 \$26460 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $762 r0 *1 579.805,864.29 sg13_lv_nmos
M$762 VSS \$26920 \$26951 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $763 r0 *1 580.655,864.195 sg13_lv_nmos
M$763 VSS \$26427 \$26965 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $764 r0 *1 580.965,864.195 sg13_lv_nmos
M$764 \$26965 \$26951 \$26478 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $765 r0 *1 582.555,864.195 sg13_lv_nmos
M$765 VSS \$25867 \$26426 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $766 r0 *1 599.085,864.355 sg13_lv_nmos
M$766 \$26957 \$25867 \$26962 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $767 r0 *1 599.595,864.355 sg13_lv_nmos
M$767 VSS \$26921 \$26962 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $768 r0 *1 600.105,864.305 sg13_lv_nmos
M$768 VSS \$26957 \$26461 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $769 r0 *1 601.395,864.29 sg13_lv_nmos
M$769 VSS \$26921 \$26952 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $770 r0 *1 602.245,864.195 sg13_lv_nmos
M$770 VSS \$25867 \$26960 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $771 r0 *1 602.555,864.195 sg13_lv_nmos
M$771 \$26960 \$26952 \$26479 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $772 r0 *1 604.145,864.195 sg13_lv_nmos
M$772 VSS \$26427 \$26428 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $773 r0 *1 620.494,863.454 sg13_lv_nmos
M$773 VSS \$26937 \$26923 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $777 r0 *1 617.465,869.102 sg13_lv_nmos
M$777 \$26994 \$26927 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $779 r0 *1 618.495,869.102 sg13_lv_nmos
M$779 \$26994 \$26993 \$27009 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $781 r0 *1 620.494,869.122 sg13_lv_nmos
M$781 VSS \$27009 \$26995 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $785 r0 *1 623.374,869.122 sg13_lv_nmos
M$785 VSS \$26995 \$26996 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $789 r0 *1 626.254,869.122 sg13_lv_nmos
M$789 VSS \$26996 \$26997 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $793 r0 *1 629.134,869.122 sg13_lv_nmos
M$793 VSS \$26997 \$26998 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $797 r0 *1 632.714,869.122 sg13_lv_nmos
M$797 VSS \$26998 \$26999 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $801 r0 *1 636.294,869.122 sg13_lv_nmos
M$801 VSS \$26999 \$26953 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $805 r0 *1 640.44,869.102 sg13_lv_nmos
M$805 \$27000 \$26953 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $807 r0 *1 641.47,869.102 sg13_lv_nmos
M$807 \$27000 \$26998 \$27010 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $809 r0 *1 643.505,869.122 sg13_lv_nmos
M$809 VSS \$27010 \$27001 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $813 r0 *1 613.57,869.127 sg13_lv_nmos
M$813 VSS \$27008 \$26954 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $815 r0 *1 615.49,869.127 sg13_lv_nmos
M$815 VSS \$26954 \$26993 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $817 r0 *1 646.325,869.128 sg13_lv_nmos
M$817 VSS \$27001 \$25867 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $825 r0 *1 1060.995,900.99 sg13_lv_nmos
M$825 \$28334 \$28308 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $826 r0 *1 1060.995,897.48 sg13_lv_nmos
M$826 \$28306 \$28308 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $827 r0 *1 478.381,936.463 sg13_lv_nmos
M$827 \$29051 \$29052 \$30346 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $828 r0 *1 483.425,932.839 sg13_lv_nmos
M$828 VSS \$29052 \$29048 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $829 r0 *1 478.382,941.223 sg13_lv_nmos
M$829 VSS \$30344 \$29390 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $830 r0 *1 480.981,941.223 sg13_lv_nmos
M$830 VSS \$29051 \$29391 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $831 r0 *1 503.35,942.602 sg13_lv_nmos
M$831 VSS \$4796 \$29392 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $832 r0 *1 504.605,942.422 sg13_lv_nmos
M$832 \$29406 \$29460 \$29418 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $833 r0 *1 504.915,942.422 sg13_lv_nmos
M$833 \$29418 \$29392 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $834 r0 *1 505.495,942.807 sg13_lv_nmos
M$834 VSS \$29430 \$29407 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $835 r0 *1 506.585,942.487 sg13_lv_nmos
M$835 VSS \$29392 \$29417 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $836 r0 *1 506.895,942.487 sg13_lv_nmos
M$836 \$29417 \$29407 \$29408 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $837 r0 *1 509.44,942.687 sg13_lv_nmos
M$837 VSS \$29409 \$29461 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $838 r0 *1 510.54,942.687 sg13_lv_nmos
M$838 VSS \$29052 \$29409 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $839 r0 *1 511.75,942.807 sg13_lv_nmos
M$839 \$29431 \$29409 \$29410 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $840 r0 *1 512.285,942.647 sg13_lv_nmos
M$840 \$29407 \$29461 \$29431 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $841 r0 *1 513.335,942.422 sg13_lv_nmos
M$841 \$29410 \$29411 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $842 r0 *1 513.845,942.422 sg13_lv_nmos
M$842 VSS \$29392 \$29420 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $843 r0 *1 514.155,942.422 sg13_lv_nmos
M$843 \$29420 \$29431 \$29411 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $844 r0 *1 516.195,942.532 sg13_lv_nmos
M$844 VSS \$29431 \$29413 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $845 r0 *1 515.175,942.582 sg13_lv_nmos
M$845 VSS \$29431 \$29412 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $847 r0 *1 517.215,942.582 sg13_lv_nmos
M$847 VSS \$29413 \$29414 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $849 r0 *1 441.615,944.16 sg13_lv_nmos
M$849 VSS \$29396 \$29397 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $853 r0 *1 444.495,944.16 sg13_lv_nmos
M$853 VSS \$29397 \$29398 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $857 r0 *1 447.375,944.16 sg13_lv_nmos
M$857 VSS \$29398 \$29399 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $861 r0 *1 450.255,944.16 sg13_lv_nmos
M$861 VSS \$29399 \$29400 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $865 r0 *1 453.135,944.16 sg13_lv_nmos
M$865 VSS \$29400 \$29401 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $869 r0 *1 456.015,944.16 sg13_lv_nmos
M$869 VSS \$29401 \$29402 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $873 r0 *1 461.775,944.16 sg13_lv_nmos
M$873 VSS \$29403 \$29404 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $877 r0 *1 464.595,944.16 sg13_lv_nmos
M$877 VSS \$29404 \$29405 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $885 r0 *1 478.179,943.829 sg13_lv_nmos
M$885 \$29424 \$29458 \$29485 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $886 r0 *1 478.381,942.756 sg13_lv_nmos
M$886 \$29390 \$29405 \$29424 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $887 r0 *1 480.981,942.752 sg13_lv_nmos
M$887 \$29391 \$29405 \$29425 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $888 r0 *1 480.985,943.845 sg13_lv_nmos
M$888 \$29425 \$29485 \$29458 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $889 r0 *1 488.224,943.679 sg13_lv_nmos
M$889 \$29426 \$29460 \$29459 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $890 r0 *1 488.24,942.636 sg13_lv_nmos
M$890 VSS \$29458 \$29426 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $891 r0 *1 491.052,942.61 sg13_lv_nmos
M$891 VSS \$29485 \$29427 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $892 r0 *1 491.053,943.68 sg13_lv_nmos
M$892 \$29427 \$29459 \$29460 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $893 r0 *1 497.502,943.659 sg13_lv_nmos
M$893 VSS \$29460 \$29428 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $894 r0 *1 498.012,943.609 sg13_lv_nmos
M$894 VSS \$29428 \$29429 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $896 r0 *1 507.67,943.212 sg13_lv_nmos
M$896 \$29406 \$29409 \$29430 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $897 r0 *1 508.18,943.212 sg13_lv_nmos
M$897 \$29430 \$29461 \$29408 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $898 r0 *1 434.915,946.5 sg13_lv_nmos
M$898 VSS \$29531 \$29423 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $900 r0 *1 436.835,946.5 sg13_lv_nmos
M$900 VSS \$29423 \$29492 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $902 r0 *1 438.7,944.185 sg13_lv_nmos
M$902 \$29456 \$29422 \$29396 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $904 r0 *1 439.73,944.185 sg13_lv_nmos
M$904 \$29456 \$29423 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $906 r0 *1 438.7,946.475 sg13_lv_nmos
M$906 \$29493 \$29492 \$29509 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $908 r0 *1 439.73,946.475 sg13_lv_nmos
M$908 \$29493 \$29402 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $910 r0 *1 441.615,946.5 sg13_lv_nmos
M$910 VSS \$29509 \$29494 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $914 r0 *1 444.495,946.5 sg13_lv_nmos
M$914 VSS \$29494 \$29495 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $918 r0 *1 447.375,946.5 sg13_lv_nmos
M$918 VSS \$29495 \$29496 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $922 r0 *1 450.255,946.5 sg13_lv_nmos
M$922 VSS \$29496 \$29497 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $926 r0 *1 453.135,946.5 sg13_lv_nmos
M$926 VSS \$29497 \$29498 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $930 r0 *1 456.015,946.5 sg13_lv_nmos
M$930 VSS \$29498 \$29422 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $934 r0 *1 458.97,944.185 sg13_lv_nmos
M$934 \$29457 \$29402 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $936 r0 *1 460,944.185 sg13_lv_nmos
M$936 \$29457 \$29400 \$29403 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $938 r0 *1 458.97,946.475 sg13_lv_nmos
M$938 \$29499 \$29422 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $940 r0 *1 460,946.475 sg13_lv_nmos
M$940 \$29499 \$29497 \$29510 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $942 r0 *1 461.775,946.5 sg13_lv_nmos
M$942 VSS \$29510 \$29500 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $946 r0 *1 464.595,946.5 sg13_lv_nmos
M$946 VSS \$29500 \$29052 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $954 r0 *1 515.91,947.59 sg13_lv_nmos
M$954 VSS \$29414 \$31708 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $956 r0 *1 436.37,962.297 sg13_lv_nmos
M$956 VSS \$29052 \$30349 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $957 r0 *1 437.455,962.397 sg13_lv_nmos
M$957 VSS \$29414 \$30350 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $958 r0 *1 438.305,962.302 sg13_lv_nmos
M$958 VSS \$29405 \$30365 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $959 r0 *1 438.615,962.302 sg13_lv_nmos
M$959 \$30365 \$30350 \$30351 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $960 r0 *1 439.93,962.467 sg13_lv_nmos
M$960 \$30352 \$29405 \$30366 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $961 r0 *1 440.44,962.467 sg13_lv_nmos
M$961 VSS \$29414 \$30366 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $962 r0 *1 440.95,962.417 sg13_lv_nmos
M$962 VSS \$30352 \$30353 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $963 r0 *1 453.856,962.757 sg13_lv_nmos
M$963 \$30340 \$29498 \$30354 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $964 r0 *1 454.365,962.757 sg13_lv_nmos
M$964 \$30354 \$29405 \$30341 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $965 r0 *1 458.256,962.737 sg13_lv_nmos
M$965 \$30342 \$29052 \$30341 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $966 r0 *1 458.765,962.737 sg13_lv_nmos
M$966 \$30341 \$4796 \$30343 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $967 r0 *1 465.452,962.297 sg13_lv_nmos
M$967 VSS \$29405 \$30355 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $968 r0 *1 466.537,962.397 sg13_lv_nmos
M$968 VSS \$29429 \$30356 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $969 r0 *1 467.387,962.302 sg13_lv_nmos
M$969 VSS \$29052 \$30369 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $970 r0 *1 467.697,962.302 sg13_lv_nmos
M$970 \$30369 \$30356 \$30357 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $971 r0 *1 469.012,962.467 sg13_lv_nmos
M$971 \$30358 \$29052 \$30371 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $972 r0 *1 469.522,962.467 sg13_lv_nmos
M$972 VSS \$29429 \$30371 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $973 r0 *1 470.032,962.417 sg13_lv_nmos
M$973 VSS \$30358 \$30359 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $974 r0 *1 482.938,962.757 sg13_lv_nmos
M$974 \$30344 \$29401 \$30360 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $975 r0 *1 483.447,962.757 sg13_lv_nmos
M$975 \$30360 \$29052 \$30361 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $976 r0 *1 487.338,962.737 sg13_lv_nmos
M$976 \$30345 \$29405 \$30361 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $977 r0 *1 487.847,962.737 sg13_lv_nmos
M$977 \$30361 \$4796 \$30346 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $978 r0 *1 445.759,966.03 sg13_lv_nmos
M$978 PAD|VLO \$30353 \$30389 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $979 r0 *1 448.177,966.092 sg13_lv_nmos
M$979 \$30389 \$29052 CORE$12 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $980 r0 *1 454.2,965.647 sg13_lv_nmos
M$980 VSS \$30340 \$30340 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $981 r0 *1 458.575,965.632 sg13_lv_nmos
M$981 VSS \$30342 \$30343 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $982 r0 *1 474.841,966.03 sg13_lv_nmos
M$982 PAD|VLO \$30359 \$30390 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $983 r0 *1 477.259,966.092 sg13_lv_nmos
M$983 \$30390 \$29405 \$30343 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $984 r0 *1 483.282,965.647 sg13_lv_nmos
M$984 VSS \$30344 \$30344 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $985 r0 *1 487.657,965.632 sg13_lv_nmos
M$985 VSS \$30345 \$30346 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $986 r0 *1 1060.995,1000.99 sg13_lv_nmos
M$986 \$31734 \$31708 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $987 r0 *1 1060.995,997.48 sg13_lv_nmos
M$987 \$31706 \$31708 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $988 r0 *1 700.255,1060.995 sg13_lv_nmos
M$988 \$16829 \$32558 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $989 r0 *1 800.255,1060.995 sg13_lv_nmos
M$989 \$27008 \$32559 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $990 r0 *1 900.255,1060.995 sg13_lv_nmos
M$990 \$29531 \$32560 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $991 r0 *1 501.765,239.055 sg13_hv_nmos
M$991 VSS CORE \$4801 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $992 r0 *1 701.765,239.055 sg13_hv_nmos
M$992 VSS CORE$1 \$4802 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $993 r0 *1 801.765,239.055 sg13_hv_nmos
M$993 VSS CORE$2 \$4803 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $994 r0 *1 901.765,239.055 sg13_hv_nmos
M$994 VSS CORE$3 \$4804 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $995 r0 *1 90.95,285.52 sg13_hv_nmos
M$995 VSS \$5434 IN6|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1015 r0 *1 1209.05,294.58 sg13_hv_nmos
M$1015 VSS \$5927 OUT6 VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999999
* device instance $1023 r0 *1 1064.68,297.64 sg13_hv_nmos
M$1023 \$5742 dout VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1024 r0 *1 1064.68,298.47 sg13_hv_nmos
M$1024 VSS \$5741 \$5752 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1025 r0 *1 1064.68,299.81 sg13_hv_nmos
M$1025 VSS \$5752 \$5927 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1026 r0 *1 1064.68,301.15 sg13_hv_nmos
M$1026 \$5947 dout VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1027 r0 *1 1064.68,301.98 sg13_hv_nmos
M$1027 VSS \$5946 \$6134 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1028 r0 *1 1064.68,303.32 sg13_hv_nmos
M$1028 VSS \$6134 \$5194 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1029 r0 *1 90.95,385.52 sg13_hv_nmos
M$1029 VSS \$9160 IN5|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1049 r0 *1 1209.05,394.58 sg13_hv_nmos
M$1049 VSS \$10159 OUT5 VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999999
* device instance $1057 r0 *1 1064.68,397.64 sg13_hv_nmos
M$1057 \$9651 \$9659 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1058 r0 *1 1064.68,398.47 sg13_hv_nmos
M$1058 VSS \$9650 \$9849 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1059 r0 *1 1064.68,399.81 sg13_hv_nmos
M$1059 VSS \$9849 \$10159 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1060 r0 *1 1064.68,401.15 sg13_hv_nmos
M$1060 \$10175 \$9659 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1061 r0 *1 1064.68,401.98 sg13_hv_nmos
M$1061 VSS \$10174 \$10185 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1062 r0 *1 1064.68,403.32 sg13_hv_nmos
M$1062 VSS \$10185 \$9150 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1063 r0 *1 90.95,485.52 sg13_hv_nmos
M$1063 VSS \$13296 IN4|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1083 r0 *1 1209.05,494.58 sg13_hv_nmos
M$1083 VSS \$13971 OUT4 VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999999
* device instance $1091 r0 *1 1064.68,497.64 sg13_hv_nmos
M$1091 \$13603 \$13736 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1092 r0 *1 1064.68,498.47 sg13_hv_nmos
M$1092 VSS \$13602 \$13787 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1093 r0 *1 1064.68,499.81 sg13_hv_nmos
M$1093 VSS \$13787 \$13971 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1094 r0 *1 1064.68,501.15 sg13_hv_nmos
M$1094 \$13983 \$13736 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1095 r0 *1 1064.68,501.98 sg13_hv_nmos
M$1095 VSS \$13982 \$13990 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1096 r0 *1 1064.68,503.32 sg13_hv_nmos
M$1096 VSS \$13990 \$13286 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1097 r0 *1 90.95,585.52 sg13_hv_nmos
M$1097 VSS \$16711 PAD|VLO VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1117 r0 *1 1139.21,663.22 sg13_hv_nmos
M$1117 VSS \$19262 \$19407 VSS sg13_hv_nmos W=108.0 L=0.5
* device instance $1123 r0 *1 1139.21,673 sg13_hv_nmos
M$1123 VSS \$19262 VSS VSS sg13_hv_nmos W=126.0 L=9.5
* device instance $1143 r0 *1 1194.53,668.155 sg13_hv_nmos
M$1143 VSS \$19407 IOVDD VSS sg13_hv_nmos W=756.7999999999977
+ L=0.5999999999999999
* device instance $1315 r0 *1 90.95,685.52 sg13_hv_nmos
M$1315 VSS \$19877 PAD|VHI VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1335 r0 *1 90.95,785.52 sg13_hv_nmos
M$1335 VSS \$23952 IN3|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1355 r0 *1 1209.05,794.58 sg13_hv_nmos
M$1355 VSS \$24435 OUT3 VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999999
* device instance $1363 r0 *1 1064.68,797.64 sg13_hv_nmos
M$1363 \$24420 \$17418 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1364 r0 *1 1064.68,798.47 sg13_hv_nmos
M$1364 VSS \$24419 \$24429 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1365 r0 *1 1064.68,799.81 sg13_hv_nmos
M$1365 VSS \$24429 \$24435 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1366 r0 *1 1064.68,801.15 sg13_hv_nmos
M$1366 \$24447 \$17418 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1367 r0 *1 1064.68,801.98 sg13_hv_nmos
M$1367 VSS \$24446 \$24454 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1368 r0 *1 1064.68,803.32 sg13_hv_nmos
M$1368 VSS \$24454 \$23485 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1369 r0 *1 510.665,859.567 sg13_hv_nmos
M$1369 \$26529 \$26529 VSS VSS sg13_hv_nmos W=33.0 L=0.9
* device instance $1377 r0 *1 530.16,859.567 sg13_hv_nmos
M$1377 \$26531 \$26529 VSS VSS sg13_hv_nmos W=33.0 L=0.9
* device instance $1385 r0 *1 495.305,859.662 sg13_hv_nmos
M$1385 \$26530 \$26529 VSS VSS sg13_hv_nmos W=33.0 L=0.9
* device instance $1393 r0 *1 506.045,858.145 sg13_hv_nmos
M$1393 VSS \$26530 \$26978 VSS sg13_hv_nmos W=1.0 L=0.44999999999999996
* device instance $1394 r0 *1 495.305,870.8 sg13_hv_nmos
M$1394 \$26955 \$26529 \$26978 VSS sg13_hv_nmos W=178.00000000000006
+ L=0.8999999999999999
* device instance $1414 r0 *1 540.27,863.82 sg13_hv_nmos
M$1414 \$25328 CORE$10 \$26531 VSS sg13_hv_nmos W=136.5 L=0.9
* device instance $1428 r0 *1 90.95,885.52 sg13_hv_nmos
M$1428 VSS \$27864 IN2|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1448 r0 *1 529.04,863.82 sg13_hv_nmos
M$1448 \$26919 PAD|VLDO \$26531 VSS sg13_hv_nmos W=136.5 L=0.9
* device instance $1462 r0 *1 1064.68,897.64 sg13_hv_nmos
M$1462 \$28307 \$28308 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1463 r0 *1 1064.68,898.47 sg13_hv_nmos
M$1463 VSS \$28306 \$28320 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1464 r0 *1 1209.05,894.58 sg13_hv_nmos
M$1464 VSS \$28323 OUT2 VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999999
* device instance $1472 r0 *1 1064.68,899.81 sg13_hv_nmos
M$1472 VSS \$28320 \$28323 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1473 r0 *1 1064.68,901.15 sg13_hv_nmos
M$1473 \$28335 \$28308 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1474 r0 *1 1064.68,901.98 sg13_hv_nmos
M$1474 VSS \$28334 \$28342 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1475 r0 *1 1064.68,903.32 sg13_hv_nmos
M$1475 VSS \$28342 \$27432 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1476 r0 *1 90.95,985.52 sg13_hv_nmos
M$1476 VSS \$31320 IN1|PAD VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $1496 r0 *1 1209.05,994.58 sg13_hv_nmos
M$1496 VSS \$31723 OUT1 VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999999
* device instance $1504 r0 *1 1064.68,997.64 sg13_hv_nmos
M$1504 \$31707 \$31708 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1505 r0 *1 1064.68,998.47 sg13_hv_nmos
M$1505 VSS \$31706 \$31717 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1506 r0 *1 1064.68,999.81 sg13_hv_nmos
M$1506 VSS \$31717 \$31723 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1507 r0 *1 1064.68,1001.15 sg13_hv_nmos
M$1507 \$31735 \$31708 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1508 r0 *1 1064.68,1001.98 sg13_hv_nmos
M$1508 VSS \$31734 \$31742 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1509 r0 *1 1064.68,1003.32 sg13_hv_nmos
M$1509 VSS \$31742 \$30871 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1510 r0 *1 701.765,1060.945 sg13_hv_nmos
M$1510 VSS CORE$13 \$32558 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $1511 r0 *1 801.765,1060.945 sg13_hv_nmos
M$1511 VSS CORE$14 \$32559 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $1512 r0 *1 901.765,1060.945 sg13_hv_nmos
M$1512 VSS CORE$15 \$32560 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $1513 r0 *1 263.22,1139.21 sg13_hv_nmos
M$1513 VSS \$33694 \$33299 VSS sg13_hv_nmos W=108.0 L=0.5
* device instance $1519 r0 *1 273,1139.21 sg13_hv_nmos
M$1519 VSS \$33694 VSS VSS sg13_hv_nmos W=126.0 L=9.5
* device instance $1526 r0 *1 563.22,1139.21 sg13_hv_nmos
M$1526 VSS \$33695 \$33300 VSS sg13_hv_nmos W=108.0 L=0.5
* device instance $1532 r0 *1 573,1139.21 sg13_hv_nmos
M$1532 VSS \$33695 VSS VSS sg13_hv_nmos W=126.0 L=9.5
* device instance $1539 r0 *1 963.22,1139.21 sg13_hv_nmos
M$1539 VSS \$33696 \$33301 VSS sg13_hv_nmos W=108.0 L=0.5
* device instance $1545 r0 *1 973,1139.21 sg13_hv_nmos
M$1545 VSS \$33696 VSS VSS sg13_hv_nmos W=126.0 L=9.5
* device instance $1591 r0 *1 268.155,1194.53 sg13_hv_nmos
M$1591 VSS \$33299 AVDD VSS sg13_hv_nmos W=756.7999999999977
+ L=0.5999999999999999
* device instance $1634 r0 *1 568.155,1194.53 sg13_hv_nmos
M$1634 VSS \$33300 IOVDD VSS sg13_hv_nmos W=756.7999999999977
+ L=0.5999999999999999
* device instance $1677 r0 *1 968.155,1194.53 sg13_hv_nmos
M$1677 VSS \$33301 VDD VSS sg13_hv_nmos W=756.7999999999977 L=0.5999999999999999
* device instance $2021 r0 *1 385.52,1209.05 sg13_hv_nmos
M$2021 VSS \$34430 PAD|VREF VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $2041 r0 *1 485.52,1209.05 sg13_hv_nmos
M$2041 VSS \$34431 PAD|VLDO VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999999
* device instance $2147 r0 *1 500.255,243.995 sg13_lv_pmos
M$2147 \$4796 \$4801 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2148 r0 *1 700.255,243.995 sg13_lv_pmos
M$2148 \$4797 \$4802 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2149 r0 *1 800.255,243.995 sg13_lv_pmos
M$2149 \$4798 \$4803 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2150 r0 *1 900.255,243.995 sg13_lv_pmos
M$2150 \$4799 \$4804 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2151 r0 *1 1056.005,297.48 sg13_lv_pmos
M$2151 \$5741 dout VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2152 r0 *1 431.875,302.8 sg13_lv_pmos
M$2152 VDD \$6129 \$6116 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2154 r0 *1 432.905,302.8 sg13_lv_pmos
M$2154 VDD \$6407 \$6116 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2156 r0 *1 434.755,302.8 sg13_lv_pmos
M$2156 VDD \$6130 \$5941 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2158 r0 *1 435.785,302.8 sg13_lv_pmos
M$2158 VDD \$6170 \$5941 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2160 r0 *1 437.56,302.8 sg13_lv_pmos
M$2160 VDD \$6116 \$5942 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2164 r0 *1 440.44,302.8 sg13_lv_pmos
M$2164 VDD \$5941 \$5943 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2168 r0 *1 443.26,302.8 sg13_lv_pmos
M$2168 VDD \$5942 \$5944 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2176 r0 *1 448.06,302.8 sg13_lv_pmos
M$2176 VDD \$5943 \$5945 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2184 r0 *1 1056.005,300.99 sg13_lv_pmos
M$2184 \$5946 dout VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2185 r0 *1 431.075,307.485 sg13_lv_pmos
M$2185 VDD \$4799 \$6165 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2187 r0 *1 433.06,307.485 sg13_lv_pmos
M$2187 VDD \$6165 \$6178 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2189 r0 *1 434.09,307.485 sg13_lv_pmos
M$2189 VDD \$6129 \$6178 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2191 r0 *1 435.865,307.485 sg13_lv_pmos
M$2191 VDD \$6178 \$6167 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2195 r0 *1 438.745,307.485 sg13_lv_pmos
M$2195 VDD \$6167 \$6168 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2199 r0 *1 441.625,307.485 sg13_lv_pmos
M$2199 VDD \$6168 \$6169 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2203 r0 *1 444.505,307.485 sg13_lv_pmos
M$2203 VDD \$6169 \$6170 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2207 r0 *1 447.385,307.485 sg13_lv_pmos
M$2207 VDD \$6170 \$6171 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2211 r0 *1 450.265,307.485 sg13_lv_pmos
M$2211 VDD \$6171 \$6130 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2215 r0 *1 456.8,304.885 sg13_lv_pmos
M$2215 VDD \$5945 \$6138 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2216 r0 *1 457.97,305.01 sg13_lv_pmos
M$2216 VDD \$5944 \$6142 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2217 r0 *1 458.48,305.01 sg13_lv_pmos
M$2217 VDD \$5926 \$6142 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2218 r0 *1 458.99,304.87 sg13_lv_pmos
M$2218 VDD \$6142 \$6139 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2219 r0 *1 460.28,304.73 sg13_lv_pmos
M$2219 \$6143 \$5926 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2220 r0 *1 460.82,304.87 sg13_lv_pmos
M$2220 VDD \$5944 \$6140 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2221 r0 *1 461.33,304.87 sg13_lv_pmos
M$2221 \$6140 \$6143 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2222 r0 *1 431.04,312.125 sg13_lv_pmos
M$2222 VDD \$6165 \$6402 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2224 r0 *1 433.025,312.125 sg13_lv_pmos
M$2224 VDD \$6130 \$6403 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2226 r0 *1 434.055,312.125 sg13_lv_pmos
M$2226 VDD \$6402 \$6403 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2228 r0 *1 435.83,312.135 sg13_lv_pmos
M$2228 VDD \$6403 \$6404 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2232 r0 *1 438.71,312.135 sg13_lv_pmos
M$2232 VDD \$6404 \$6405 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2236 r0 *1 441.59,312.135 sg13_lv_pmos
M$2236 VDD \$6405 \$6406 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2240 r0 *1 444.47,312.135 sg13_lv_pmos
M$2240 VDD \$6406 \$6407 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2244 r0 *1 447.35,312.135 sg13_lv_pmos
M$2244 VDD \$6407 \$6408 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2248 r0 *1 450.23,312.135 sg13_lv_pmos
M$2248 VDD \$6408 \$6129 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2252 r0 *1 457.62,310.765 sg13_lv_pmos
M$2252 \$6193 \$6140 PAD|VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2253 r0 *1 460.105,309.515 sg13_lv_pmos
M$2253 \$6193 \$6138 \$6197 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2256 r0 *1 431.695,323.31 sg13_lv_pmos
M$2256 VDD \$5944 \$6971 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2257 r0 *1 432.865,323.435 sg13_lv_pmos
M$2257 VDD \$5945 \$6972 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2258 r0 *1 433.375,323.435 sg13_lv_pmos
M$2258 VDD \$6782 \$6972 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2259 r0 *1 433.885,323.295 sg13_lv_pmos
M$2259 VDD \$6972 \$6973 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2260 r0 *1 435.175,323.155 sg13_lv_pmos
M$2260 \$6974 \$6782 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2261 r0 *1 435.715,323.295 sg13_lv_pmos
M$2261 VDD \$5945 \$6975 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2262 r0 *1 436.225,323.295 sg13_lv_pmos
M$2262 \$6975 \$6974 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2263 r0 *1 451.11,327.385 sg13_lv_pmos
M$2263 VDD \$5944 \$7301 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2264 r0 *1 452.55,327.385 sg13_lv_pmos
M$2264 VDD \$4796 \$7302 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2265 r0 *1 454.96,327.385 sg13_lv_pmos
M$2265 VDD \$7385 \$7322 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2266 r0 *1 453.94,327.37 sg13_lv_pmos
M$2266 VDD \$7322 \$5926 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2268 r0 *1 461.43,327.36 sg13_lv_pmos
M$2268 \$7339 \$7305 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2269 r0 *1 462.155,327.36 sg13_lv_pmos
M$2269 VDD \$5944 \$7305 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2270 r0 *1 465.395,311.56 sg13_lv_pmos
M$2270 AVDD \$6144 \$6144 AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2274 r0 *1 469.615,311.56 sg13_lv_pmos
M$2274 AVDD \$6118 \$6117 AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2278 r0 *1 468.43,327.37 sg13_lv_pmos
M$2278 VDD \$7309 \$6782 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2280 r0 *1 470.55,327.37 sg13_lv_pmos
M$2280 VDD \$6782 dout VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2282 r0 *1 435,327.94 sg13_lv_pmos
M$2282 \$7314 \$6971 CORE$4 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2285 r0 *1 456.085,327.12 sg13_lv_pmos
M$2285 VDD \$7385 \$7303 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2286 r0 *1 456.595,327.12 sg13_lv_pmos
M$2286 VDD \$7302 \$7303 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2287 r0 *1 457.045,327.41 sg13_lv_pmos
M$2287 VDD \$7323 \$7304 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2288 r0 *1 458.095,327.485 sg13_lv_pmos
M$2288 \$7323 \$7302 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2289 r0 *1 458.83,327.485 sg13_lv_pmos
M$2289 VDD \$7304 \$7349 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2290 r0 *1 459.22,327.485 sg13_lv_pmos
M$2290 \$7349 \$7305 \$7323 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2291 r0 *1 459.73,327.485 sg13_lv_pmos
M$2291 \$7323 \$7339 \$7303 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2292 r0 *1 464.285,327.105 sg13_lv_pmos
M$2292 \$7316 \$7339 \$7352 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2293 r0 *1 464.665,327.105 sg13_lv_pmos
M$2293 \$7352 \$7307 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2294 r0 *1 465.275,327.105 sg13_lv_pmos
M$2294 VDD \$7302 \$7307 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2295 r0 *1 465.785,327.105 sg13_lv_pmos
M$2295 VDD \$7316 \$7307 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2296 r0 *1 467.345,327.21 sg13_lv_pmos
M$2296 VDD \$7316 \$7309 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2297 r0 *1 466.325,327.27 sg13_lv_pmos
M$2297 VDD \$7316 \$7308 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2299 r0 *1 463.59,327.395 sg13_lv_pmos
M$2299 \$7304 \$7305 \$7316 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2300 r0 *1 432.515,329.19 sg13_lv_pmos
M$2300 \$7314 \$6975 PAD|VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2301 r0 *1 440.29,329.985 sg13_lv_pmos
M$2301 AVDD \$7039 \$7039 AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2305 r0 *1 460.335,334.2 sg13_lv_pmos
M$2305 AVDD \$5945 \$7383 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2306 r0 *1 460.845,334.2 sg13_lv_pmos
M$2306 \$7383 \$7378 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2307 r0 *1 463.38,334.225 sg13_lv_pmos
M$2307 AVDD \$7383 \$7378 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2308 r0 *1 463.89,334.225 sg13_lv_pmos
M$2308 \$7378 \$5945 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2309 r0 *1 467.145,334.24 sg13_lv_pmos
M$2309 VDD \$7378 \$7384 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2310 r0 *1 467.655,334.24 sg13_lv_pmos
M$2310 \$7384 \$7385 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2311 r0 *1 470.18,334.24 sg13_lv_pmos
M$2311 VDD \$7384 \$7385 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2312 r0 *1 470.69,334.24 sg13_lv_pmos
M$2312 \$7385 \$7383 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2313 r0 *1 444.51,329.985 sg13_lv_pmos
M$2313 AVDD \$6783 \$6197 AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2317 r0 *1 458.31,333.385 sg13_lv_pmos
M$2317 \$7364 \$7301 \$6117 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2320 r0 *1 464.231,395.258 sg13_lv_pmos
M$2320 \$9628 \$9632 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2321 r0 *1 464.741,395.398 sg13_lv_pmos
M$2321 VDD \$9659 \$9632 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2322 r0 *1 465.251,395.398 sg13_lv_pmos
M$2322 \$9632 \$10180 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2323 r0 *1 476.371,395.398 sg13_lv_pmos
M$2323 VDD \$9658 \$9633 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2324 r0 *1 476.881,395.398 sg13_lv_pmos
M$2324 VDD \$9635 \$9633 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2325 r0 *1 477.391,395.258 sg13_lv_pmos
M$2325 VDD \$9633 \$9629 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2326 r0 *1 463.96,399.379 sg13_lv_pmos
M$2326 \$9634 \$9842 CORE$5 AVDD sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2330 r0 *1 476.132,399.379 sg13_lv_pmos
M$2330 \$9848 \$9843 \$10410 AVDD sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2334 r0 *1 1056.005,397.48 sg13_lv_pmos
M$2334 \$9650 \$9659 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2335 r0 *1 1056.005,400.99 sg13_lv_pmos
M$2335 \$10174 \$9659 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2336 r0 *1 466.182,407.008 sg13_lv_pmos
M$2336 PAD|VHI \$10206 \$9634 AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2337 r0 *1 475.44,407.008 sg13_lv_pmos
M$2337 \$9848 \$10207 PAD|VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2338 r0 *1 462.071,407.38 sg13_lv_pmos
M$2338 \$10208 \$9659 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2339 r0 *1 462.611,407.52 sg13_lv_pmos
M$2339 VDD \$10180 \$10206 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2340 r0 *1 463.121,407.52 sg13_lv_pmos
M$2340 \$10206 \$10208 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2341 r0 *1 479.551,407.38 sg13_lv_pmos
M$2341 VDD \$9635 \$10209 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2342 r0 *1 478.501,407.52 sg13_lv_pmos
M$2342 VDD \$10209 \$10207 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2343 r0 *1 479.011,407.52 sg13_lv_pmos
M$2343 \$10207 \$9658 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2344 r0 *1 441.983,411.264 sg13_lv_pmos
M$2344 \$10183 \$10183 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2348 r0 *1 458.733,407.535 sg13_lv_pmos
M$2348 VDD \$9658 \$9842 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2349 r0 *1 482.889,407.535 sg13_lv_pmos
M$2349 \$9843 \$10180 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2350 r0 *1 493.999,411.264 sg13_lv_pmos
M$2350 \$10184 \$10184 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2354 r0 *1 441.983,420.81 sg13_lv_pmos
M$2354 \$10410 \$9622 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2358 r0 *1 493.999,420.81 sg13_lv_pmos
M$2358 \$10411 \$9625 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2362 r0 *1 452.732,432.655 sg13_lv_pmos
M$2362 VDD \$11326 \$10926 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2364 r0 *1 453.762,432.655 sg13_lv_pmos
M$2364 VDD \$11335 \$10926 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2366 r0 *1 455.996,432.655 sg13_lv_pmos
M$2366 VDD \$10926 \$10927 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2370 r0 *1 459.411,432.655 sg13_lv_pmos
M$2370 VDD \$10927 \$10928 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2374 r0 *1 462.647,432.655 sg13_lv_pmos
M$2374 VDD \$10928 \$10929 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2378 r0 *1 466.172,432.655 sg13_lv_pmos
M$2378 VDD \$10929 \$10930 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2382 r0 *1 470.029,432.655 sg13_lv_pmos
M$2382 VDD \$10930 \$10931 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2386 r0 *1 473.998,432.655 sg13_lv_pmos
M$2386 VDD \$10931 \$10932 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2390 r0 *1 477.918,432.655 sg13_lv_pmos
M$2390 VDD \$10932 \$10934 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2392 r0 *1 478.948,432.655 sg13_lv_pmos
M$2392 VDD \$10930 \$10934 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2394 r0 *1 481.602,432.655 sg13_lv_pmos
M$2394 VDD \$10934 \$10935 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2398 r0 *1 484.998,432.655 sg13_lv_pmos
M$2398 VDD \$10935 \$10180 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2406 r0 *1 446.833,440.623 sg13_lv_pmos
M$2406 VDD \$4798 \$11326 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2408 r0 *1 449.354,440.623 sg13_lv_pmos
M$2408 VDD \$11326 \$11327 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2410 r0 *1 452.01,440.623 sg13_lv_pmos
M$2410 VDD \$11327 \$11329 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2412 r0 *1 453.04,440.623 sg13_lv_pmos
M$2412 VDD \$10932 \$11329 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2414 r0 *1 455.373,440.624 sg13_lv_pmos
M$2414 VDD \$11329 \$11330 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2418 r0 *1 459.841,440.624 sg13_lv_pmos
M$2418 VDD \$11330 \$11331 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2422 r0 *1 463.257,440.624 sg13_lv_pmos
M$2422 VDD \$11331 \$11332 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2426 r0 *1 466.777,440.624 sg13_lv_pmos
M$2426 VDD \$11332 \$11333 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2430 r0 *1 470.634,440.624 sg13_lv_pmos
M$2430 VDD \$11333 \$11334 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2434 r0 *1 474.603,440.624 sg13_lv_pmos
M$2434 VDD \$11334 \$11335 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2438 r0 *1 478.273,440.624 sg13_lv_pmos
M$2438 VDD \$11335 \$11337 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2440 r0 *1 479.303,440.624 sg13_lv_pmos
M$2440 VDD \$11333 \$11337 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2442 r0 *1 481.957,440.624 sg13_lv_pmos
M$2442 VDD \$11337 \$11338 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2446 r0 *1 485.353,440.624 sg13_lv_pmos
M$2446 VDD \$11338 \$9658 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2454 r0 *1 448.934,453.235 sg13_lv_pmos
M$2454 \$11717 \$11690 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2455 r0 *1 448.934,459.035 sg13_lv_pmos
M$2455 \$12329 \$11646 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2456 r0 *1 450.344,448.117 sg13_lv_pmos
M$2456 VDD \$11717 \$11666 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2457 r0 *1 449.324,448.102 sg13_lv_pmos
M$2457 VDD \$11666 \$9635 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2459 r0 *1 452.214,447.852 sg13_lv_pmos
M$2459 VDD \$11717 \$11649 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2460 r0 *1 452.724,447.852 sg13_lv_pmos
M$2460 VDD \$11650 \$11649 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2461 r0 *1 453.174,448.142 sg13_lv_pmos
M$2461 VDD \$11686 \$11651 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2462 r0 *1 452.376,459.035 sg13_lv_pmos
M$2462 VDD \$11717 \$12329 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2463 r0 *1 452.376,453.235 sg13_lv_pmos
M$2463 VDD \$12329 \$11717 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2464 r0 *1 454.224,448.217 sg13_lv_pmos
M$2464 \$11686 \$11650 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2465 r0 *1 454.959,448.217 sg13_lv_pmos
M$2465 VDD \$11651 \$11692 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2466 r0 *1 455.349,448.217 sg13_lv_pmos
M$2466 \$11692 \$11653 \$11686 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2467 r0 *1 455.859,448.217 sg13_lv_pmos
M$2467 \$11686 \$11667 \$11649 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2468 r0 *1 457.559,448.092 sg13_lv_pmos
M$2468 \$11667 \$11653 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2469 r0 *1 458.284,448.092 sg13_lv_pmos
M$2469 VDD \$9658 \$11653 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2470 r0 *1 460.414,447.837 sg13_lv_pmos
M$2470 \$11668 \$11667 \$11695 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2471 r0 *1 460.794,447.837 sg13_lv_pmos
M$2471 \$11695 \$11655 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2472 r0 *1 461.404,447.837 sg13_lv_pmos
M$2472 VDD \$11650 \$11655 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2473 r0 *1 461.914,447.837 sg13_lv_pmos
M$2473 VDD \$11668 \$11655 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2474 r0 *1 463.474,447.942 sg13_lv_pmos
M$2474 VDD \$11668 \$11657 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2475 r0 *1 462.454,448.002 sg13_lv_pmos
M$2475 VDD \$11668 \$11656 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2477 r0 *1 459.719,448.127 sg13_lv_pmos
M$2477 \$11651 \$11653 \$11668 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2478 r0 *1 464.559,448.102 sg13_lv_pmos
M$2478 VDD \$11657 \$9659 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2480 r0 *1 467.715,448.117 sg13_lv_pmos
M$2480 VDD \$4796 \$11650 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2481 r0 *1 469.15,448.117 sg13_lv_pmos
M$2481 VDD \$9658 \$11658 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2482 r0 *1 470.978,449.053 sg13_lv_pmos
M$2482 \$10411 \$11658 \$11659 AVDD sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2483 r0 *1 481.568,446.364 sg13_lv_pmos
M$2483 AVDD \$11690 \$11646 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2484 r0 *1 481.568,452.025 sg13_lv_pmos
M$2484 AVDD \$11646 \$11690 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2485 r0 *1 486.915,446.364 sg13_lv_pmos
M$2485 \$11646 \$10180 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2486 r0 *1 486.915,452.025 sg13_lv_pmos
M$2486 \$11690 \$10180 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2487 r0 *1 1056.005,497.48 sg13_lv_pmos
M$2487 \$13602 \$13736 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2488 r0 *1 1056.005,500.99 sg13_lv_pmos
M$2488 \$13982 \$13736 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2489 r0 *1 484.613,506.087 sg13_lv_pmos
M$2489 VDD \$14004 \$14005 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2490 r0 *1 485.123,506.087 sg13_lv_pmos
M$2490 \$14005 \$14016 \$14006 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2491 r0 *1 485.773,506.417 sg13_lv_pmos
M$2491 \$14006 \$13999 \$14041 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2492 r0 *1 486.108,506.417 sg13_lv_pmos
M$2492 \$14041 \$14007 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2493 r0 *1 486.618,506.417 sg13_lv_pmos
M$2493 VDD \$13993 \$14007 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2494 r0 *1 487.128,506.417 sg13_lv_pmos
M$2494 VDD \$14006 \$14007 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2495 r0 *1 487.688,506.252 sg13_lv_pmos
M$2495 VDD \$14006 \$14008 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2496 r0 *1 497.628,506.266 sg13_lv_pmos
M$2496 VDD \$14233 \$14030 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2497 r0 *1 496.608,506.251 sg13_lv_pmos
M$2497 VDD \$14030 \$14011 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2499 r0 *1 489.163,506.392 sg13_lv_pmos
M$2499 VDD \$14006 \$14009 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2500 r0 *1 489.673,506.252 sg13_lv_pmos
M$2500 VDD \$14009 \$14010 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2501 r0 *1 491.888,506.252 sg13_lv_pmos
M$2501 VDD \$14010 \$13736 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2503 r0 *1 476.778,506.267 sg13_lv_pmos
M$2503 VDD \$14713 \$14002 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2504 r0 *1 480.303,506.312 sg13_lv_pmos
M$2504 \$14016 \$14713 VDD VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2505 r0 *1 480.813,506.312 sg13_lv_pmos
M$2505 VDD \$14016 \$13999 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2506 r0 *1 481.973,506.377 sg13_lv_pmos
M$2506 \$14003 \$13999 \$14004 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2507 r0 *1 482.483,506.377 sg13_lv_pmos
M$2507 \$14004 \$14016 \$14039 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2508 r0 *1 482.858,506.377 sg13_lv_pmos
M$2508 \$14039 \$14005 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2509 r0 *1 483.433,506.377 sg13_lv_pmos
M$2509 VDD \$13993 \$14004 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2510 r0 *1 494.703,506.266 sg13_lv_pmos
M$2510 VDD \$4796 \$13993 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2511 r0 *1 478.773,506.602 sg13_lv_pmos
M$2511 VDD \$14233 \$14003 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2512 r0 *1 479.283,506.602 sg13_lv_pmos
M$2512 \$14003 \$13993 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2513 r0 *1 481.401,518.61 sg13_lv_pmos
M$2513 \$14206 \$14250 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2514 r0 *1 482.801,518.61 sg13_lv_pmos
M$2514 AVDD \$14232 \$14206 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2515 r0 *1 484.201,518.61 sg13_lv_pmos
M$2515 \$14232 \$14206 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2516 r0 *1 485.601,518.61 sg13_lv_pmos
M$2516 AVDD \$14250 \$14232 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2517 r0 *1 489.122,508.991 sg13_lv_pmos
M$2517 \$14121 \$14002 \$14122 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2520 r0 *1 488.259,518.61 sg13_lv_pmos
M$2520 \$14209 \$14232 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2521 r0 *1 489.659,518.61 sg13_lv_pmos
M$2521 VDD \$14233 \$14209 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2522 r0 *1 491.059,518.61 sg13_lv_pmos
M$2522 \$14233 \$14209 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2523 r0 *1 492.459,518.61 sg13_lv_pmos
M$2523 VDD \$14206 \$14233 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2524 r0 *1 435.35,517.186 sg13_lv_pmos
M$2524 VDD \$14709 \$14241 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2526 r0 *1 436.38,517.186 sg13_lv_pmos
M$2526 VDD \$14258 \$14241 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2528 r0 *1 438.155,517.186 sg13_lv_pmos
M$2528 VDD \$14241 \$14242 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2532 r0 *1 441.035,517.186 sg13_lv_pmos
M$2532 VDD \$14242 \$14243 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2536 r0 *1 443.915,517.186 sg13_lv_pmos
M$2536 VDD \$14243 \$14244 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2540 r0 *1 446.795,517.186 sg13_lv_pmos
M$2540 VDD \$14244 \$14245 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2544 r0 *1 449.675,517.186 sg13_lv_pmos
M$2544 VDD \$14245 \$14246 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2548 r0 *1 452.555,517.186 sg13_lv_pmos
M$2548 VDD \$14246 \$14247 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2552 r0 *1 455.51,517.186 sg13_lv_pmos
M$2552 VDD \$14247 \$14248 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2554 r0 *1 456.54,517.186 sg13_lv_pmos
M$2554 VDD \$14245 \$14248 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2556 r0 *1 458.315,517.186 sg13_lv_pmos
M$2556 VDD \$14248 \$14249 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2560 r0 *1 461.135,517.186 sg13_lv_pmos
M$2560 VDD \$14249 \$14250 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2568 r0 *1 431.445,522.941 sg13_lv_pmos
M$2568 VDD \$4797 \$14258 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2570 r0 *1 432.935,536.781 sg13_lv_pmos
M$2570 \$15033 \$14010 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2571 r0 *1 433.475,536.921 sg13_lv_pmos
M$2571 VDD \$14250 \$15027 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2572 r0 *1 433.985,536.921 sg13_lv_pmos
M$2572 \$15027 \$15033 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2573 r0 *1 433.365,522.941 sg13_lv_pmos
M$2573 VDD \$14258 \$14702 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2575 r0 *1 435.35,522.941 sg13_lv_pmos
M$2575 VDD \$14247 \$14718 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2577 r0 *1 436.38,522.941 sg13_lv_pmos
M$2577 VDD \$14702 \$14718 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2579 r0 *1 438.155,522.941 sg13_lv_pmos
M$2579 VDD \$14718 \$14704 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2583 r0 *1 441.035,522.941 sg13_lv_pmos
M$2583 VDD \$14704 \$14705 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2587 r0 *1 443.915,522.941 sg13_lv_pmos
M$2587 VDD \$14705 \$14706 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2591 r0 *1 446.795,522.941 sg13_lv_pmos
M$2591 VDD \$14706 \$14707 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2595 r0 *1 449.675,522.941 sg13_lv_pmos
M$2595 VDD \$14707 \$14708 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2599 r0 *1 452.555,522.941 sg13_lv_pmos
M$2599 VDD \$14708 \$14709 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2603 r0 *1 455.51,522.941 sg13_lv_pmos
M$2603 VDD \$14709 \$14711 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2605 r0 *1 456.54,522.941 sg13_lv_pmos
M$2605 VDD \$14707 \$14711 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2607 r0 *1 458.315,522.941 sg13_lv_pmos
M$2607 VDD \$14711 \$14712 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2611 r0 *1 461.135,522.941 sg13_lv_pmos
M$2611 VDD \$14712 \$14713 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2619 r0 *1 467.935,536.781 sg13_lv_pmos
M$2619 \$15035 \$14011 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2620 r0 *1 468.475,536.921 sg13_lv_pmos
M$2620 VDD \$14713 \$15031 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2621 r0 *1 468.985,536.921 sg13_lv_pmos
M$2621 \$15031 \$15035 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2622 r0 *1 431.51,536.936 sg13_lv_pmos
M$2622 VDD \$14713 \$15026 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2623 r0 *1 435.785,537.061 sg13_lv_pmos
M$2623 VDD \$14250 \$15034 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2624 r0 *1 436.295,537.061 sg13_lv_pmos
M$2624 VDD \$14010 \$15034 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2625 r0 *1 436.805,536.921 sg13_lv_pmos
M$2625 VDD \$15034 \$15028 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2626 r0 *1 452.577,539.206 sg13_lv_pmos
M$2626 \$15048 \$15047 AVDD AVDD sg13_lv_pmos W=10.5 L=1.5
* device instance $2630 r0 *1 466.51,536.936 sg13_lv_pmos
M$2630 VDD \$14250 \$15030 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2631 r0 *1 470.785,537.061 sg13_lv_pmos
M$2631 VDD \$14713 \$15036 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2632 r0 *1 471.295,537.061 sg13_lv_pmos
M$2632 VDD \$14011 \$15036 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2633 r0 *1 471.805,536.921 sg13_lv_pmos
M$2633 VDD \$15036 \$15032 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2634 r0 *1 487.577,539.206 sg13_lv_pmos
M$2634 \$14121 \$15049 AVDD AVDD sg13_lv_pmos W=10.5 L=1.5
* device instance $2638 r0 *1 440.927,539.221 sg13_lv_pmos
M$2638 \$15029 \$15029 AVDD AVDD sg13_lv_pmos W=10.5 L=1.5
* device instance $2642 r0 *1 475.927,539.221 sg13_lv_pmos
M$2642 \$14194 \$14194 AVDD AVDD sg13_lv_pmos W=10.5 L=1.5
* device instance $2646 r0 *1 434.41,549.416 sg13_lv_pmos
M$2646 \$15336 \$15027 PAD|VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2647 r0 *1 436.765,548.916 sg13_lv_pmos
M$2647 \$15336 \$15026 CORE$6 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2650 r0 *1 469.41,549.416 sg13_lv_pmos
M$2650 \$15076 \$15031 PAD|VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2651 r0 *1 471.765,548.916 sg13_lv_pmos
M$2651 \$15076 \$15030 \$15048 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2654 r0 *1 449.83,598.84 sg13_lv_pmos
M$2654 VDD \$17062 \$16932 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2656 r0 *1 450.86,598.84 sg13_lv_pmos
M$2656 VDD \$16931 \$16932 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2658 r0 *1 452.635,598.84 sg13_lv_pmos
M$2658 VDD \$16932 \$16922 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2662 r0 *1 455.515,598.84 sg13_lv_pmos
M$2662 VDD \$16922 \$16923 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2666 r0 *1 458.395,598.84 sg13_lv_pmos
M$2666 VDD \$16923 \$16924 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2670 r0 *1 461.275,598.84 sg13_lv_pmos
M$2670 VDD \$16924 \$16925 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2674 r0 *1 464.155,598.84 sg13_lv_pmos
M$2674 VDD \$16925 \$16926 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2678 r0 *1 467.035,598.84 sg13_lv_pmos
M$2678 VDD \$16926 \$16927 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2682 r0 *1 469.99,598.84 sg13_lv_pmos
M$2682 VDD \$16927 \$16933 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2684 r0 *1 471.02,598.84 sg13_lv_pmos
M$2684 VDD \$16925 \$16933 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2686 r0 *1 472.795,598.84 sg13_lv_pmos
M$2686 VDD \$16933 \$16929 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2690 r0 *1 475.615,598.84 sg13_lv_pmos
M$2690 VDD \$16929 \$16930 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2698 r0 *1 445.925,604.64 sg13_lv_pmos
M$2698 VDD \$16829 \$16931 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2700 r0 *1 447.845,604.64 sg13_lv_pmos
M$2700 VDD \$16931 \$17055 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2702 r0 *1 449.83,604.64 sg13_lv_pmos
M$2702 VDD \$16927 \$17066 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2704 r0 *1 450.86,604.64 sg13_lv_pmos
M$2704 VDD \$17055 \$17066 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2706 r0 *1 452.635,604.64 sg13_lv_pmos
M$2706 VDD \$17066 \$17057 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2710 r0 *1 455.515,604.64 sg13_lv_pmos
M$2710 VDD \$17057 \$17058 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2714 r0 *1 458.395,604.64 sg13_lv_pmos
M$2714 VDD \$17058 \$17059 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2718 r0 *1 461.275,604.64 sg13_lv_pmos
M$2718 VDD \$17059 \$17060 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2722 r0 *1 464.155,604.64 sg13_lv_pmos
M$2722 VDD \$17060 \$17061 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2726 r0 *1 467.035,604.64 sg13_lv_pmos
M$2726 VDD \$17061 \$17062 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2730 r0 *1 469.99,604.64 sg13_lv_pmos
M$2730 VDD \$17062 \$17067 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2732 r0 *1 471.02,604.64 sg13_lv_pmos
M$2732 VDD \$17060 \$17067 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2734 r0 *1 472.795,604.64 sg13_lv_pmos
M$2734 VDD \$17067 \$17064 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2738 r0 *1 475.615,604.64 sg13_lv_pmos
M$2738 VDD \$17064 \$17065 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2746 r0 *1 433.28,618.09 sg13_lv_pmos
M$2746 VDD \$17065 \$17383 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2747 r0 *1 434.36,617.935 sg13_lv_pmos
M$2747 \$17384 \$17226 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2748 r0 *1 434.9,618.075 sg13_lv_pmos
M$2748 VDD \$16930 \$17381 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2749 r0 *1 435.41,618.075 sg13_lv_pmos
M$2749 \$17381 \$17384 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2750 r0 *1 434.995,621.675 sg13_lv_pmos
M$2750 CORE$9 \$17383 \$17495 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2753 r0 *1 436.85,618.215 sg13_lv_pmos
M$2753 VDD \$16930 \$17388 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2754 r0 *1 437.36,618.215 sg13_lv_pmos
M$2754 VDD \$17226 \$17388 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2755 r0 *1 437.87,618.075 sg13_lv_pmos
M$2755 VDD \$17388 \$17369 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2756 r0 *1 439.97,617.765 sg13_lv_pmos
M$2756 PAD|VHI \$17381 \$17495 AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2757 r0 *1 469.335,618.09 sg13_lv_pmos
M$2757 VDD \$16930 \$17385 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2758 r0 *1 470.415,617.935 sg13_lv_pmos
M$2758 \$17386 \$17355 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2759 r0 *1 470.955,618.075 sg13_lv_pmos
M$2759 VDD \$17065 \$17382 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2760 r0 *1 471.465,618.075 sg13_lv_pmos
M$2760 \$17382 \$17386 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2761 r0 *1 471.05,621.675 sg13_lv_pmos
M$2761 \$17496 \$17385 \$17540 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2764 r0 *1 472.905,618.215 sg13_lv_pmos
M$2764 VDD \$17065 \$17389 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2765 r0 *1 473.415,618.215 sg13_lv_pmos
M$2765 VDD \$17355 \$17389 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2766 r0 *1 473.925,618.075 sg13_lv_pmos
M$2766 VDD \$17389 \$17371 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2767 r0 *1 476.025,617.765 sg13_lv_pmos
M$2767 PAD|VHI \$17382 \$17540 AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2768 r0 *1 505.15,621.115 sg13_lv_pmos
M$2768 \$17662 \$17387 \$17497 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2771 r0 *1 505.435,618.205 sg13_lv_pmos
M$2771 VDD \$17065 \$17387 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2772 r0 *1 520.805,621.42 sg13_lv_pmos
M$2772 VDD \$17650 \$17541 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2773 r0 *1 521.315,621.42 sg13_lv_pmos
M$2773 VDD \$17536 \$17541 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2774 r0 *1 521.765,621.71 sg13_lv_pmos
M$2774 VDD \$17663 \$17542 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2775 r0 *1 526.15,621.66 sg13_lv_pmos
M$2775 \$17651 \$17543 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2776 r0 *1 526.875,621.66 sg13_lv_pmos
M$2776 VDD \$17065 \$17543 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2777 r0 *1 529.005,621.405 sg13_lv_pmos
M$2777 \$17652 \$17651 \$17676 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2778 r0 *1 529.385,621.405 sg13_lv_pmos
M$2778 \$17676 \$17545 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2779 r0 *1 529.995,621.405 sg13_lv_pmos
M$2779 VDD \$17536 \$17545 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2780 r0 *1 530.505,621.405 sg13_lv_pmos
M$2780 VDD \$17652 \$17545 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2781 r0 *1 532.065,621.51 sg13_lv_pmos
M$2781 VDD \$17652 \$17547 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2782 r0 *1 531.045,621.57 sg13_lv_pmos
M$2782 VDD \$17652 \$17546 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2784 r0 *1 528.31,621.695 sg13_lv_pmos
M$2784 \$17542 \$17543 \$17652 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2785 r0 *1 533.15,621.67 sg13_lv_pmos
M$2785 VDD \$17547 \$17226 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2787 r0 *1 535.2,621.67 sg13_lv_pmos
M$2787 VDD \$17226 \$17418 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2789 r0 *1 536.99,621.68 sg13_lv_pmos
M$2789 \$17536 \$4796 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2790 r0 *1 456.64,625.975 sg13_lv_pmos
M$2790 \$17496 \$17412 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2794 r0 *1 462.64,625.975 sg13_lv_pmos
M$2794 \$17370 \$17370 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2798 r0 *1 492.695,625.975 sg13_lv_pmos
M$2798 \$17497 \$17413 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2802 r0 *1 498.695,625.975 sg13_lv_pmos
M$2802 \$17372 \$17372 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $2806 r0 *1 521.51,632.615 sg13_lv_pmos
M$2806 VDD \$17900 \$17727 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2807 r0 *1 522.815,621.785 sg13_lv_pmos
M$2807 \$17663 \$17536 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2808 r0 *1 523.55,621.785 sg13_lv_pmos
M$2808 VDD \$17542 \$17684 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2809 r0 *1 523.94,621.785 sg13_lv_pmos
M$2809 \$17684 \$17543 \$17663 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2810 r0 *1 524.45,621.785 sg13_lv_pmos
M$2810 \$17663 \$17651 \$17541 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2811 r0 *1 524.18,632.615 sg13_lv_pmos
M$2811 \$17727 \$17650 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2812 r0 *1 528.19,632.615 sg13_lv_pmos
M$2812 VDD \$17727 \$17650 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2813 r0 *1 530.86,632.615 sg13_lv_pmos
M$2813 \$17650 \$17899 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2814 r0 *1 534.455,625.47 sg13_lv_pmos
M$2814 VDD \$17703 \$17355 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2816 r0 *1 534.47,626.49 sg13_lv_pmos
M$2816 VDD \$17650 \$17703 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2817 r0 *1 508.41,633.315 sg13_lv_pmos
M$2817 AVDD \$16930 \$17899 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2818 r0 *1 511.055,633.315 sg13_lv_pmos
M$2818 \$17899 \$17900 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2819 r0 *1 513.41,633.315 sg13_lv_pmos
M$2819 AVDD \$17899 \$17900 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2820 r0 *1 516.045,633.315 sg13_lv_pmos
M$2820 \$17900 \$16930 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2821 r0 *1 1056.005,797.48 sg13_lv_pmos
M$2821 \$24419 \$17418 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2822 r0 *1 1056.005,800.99 sg13_lv_pmos
M$2822 \$24446 \$17418 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2823 r0 *1 633.21,840.21 sg13_lv_pmos
M$2823 PAD|VLDO \$25483 \$25483 PAD|VLDO sg13_lv_pmos W=10.0 L=1.5
* device instance $2825 r0 *1 630.06,845.38 sg13_lv_pmos
M$2825 \$25822 \$25853 \$25487 PAD|VLDO sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2827 r0 *1 622.075,848.775 sg13_lv_pmos
M$2827 PAD|VLDO \$26427 \$25839 PAD|VLDO sg13_lv_pmos W=4.0 L=0.13
* device instance $2829 r0 *1 624.015,848.775 sg13_lv_pmos
M$2829 PAD|VLDO \$25838 \$25839 PAD|VLDO sg13_lv_pmos W=4.0 L=0.13
* device instance $2831 r0 *1 625.955,848.775 sg13_lv_pmos
M$2831 PAD|VLDO \$25839 \$25838 PAD|VLDO sg13_lv_pmos W=4.0 L=0.13
* device instance $2833 r0 *1 627.895,848.775 sg13_lv_pmos
M$2833 PAD|VLDO \$26427 \$25838 PAD|VLDO sg13_lv_pmos W=4.0 L=0.13
* device instance $2835 r0 *1 631.3,848.775 sg13_lv_pmos
M$2835 VDD \$25838 \$25850 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2837 r0 *1 633.24,848.775 sg13_lv_pmos
M$2837 VDD \$25840 \$25850 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2839 r0 *1 635.18,848.775 sg13_lv_pmos
M$2839 VDD \$25850 \$25840 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2841 r0 *1 637.12,848.775 sg13_lv_pmos
M$2841 VDD \$25839 \$25840 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2843 r0 *1 585.345,849.525 sg13_lv_pmos
M$2843 \$25848 \$26426 CORE$11 PAD|VLDO sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2845 r0 *1 586.14,853.855 sg13_lv_pmos
M$2845 PAD|VHI \$26478 \$25848 PAD|VLDO sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2846 r0 *1 592.87,850.555 sg13_lv_pmos
M$2846 PAD|VLDO \$25489 \$25833 PAD|VLDO sg13_lv_pmos W=10.0 L=1.5
* device instance $2848 r0 *1 606.935,849.525 sg13_lv_pmos
M$2848 \$25849 \$26428 \$25833 PAD|VLDO sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2850 r0 *1 607.73,853.855 sg13_lv_pmos
M$2850 PAD|VHI \$26479 \$25849 PAD|VLDO sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2851 r0 *1 614.46,850.555 sg13_lv_pmos
M$2851 PAD|VLDO \$25490 \$25822 PAD|VLDO sg13_lv_pmos W=10.0 L=1.5
* device instance $2853 r0 *1 628.87,853.995 sg13_lv_pmos
M$2853 \$26497 \$26450 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2854 r0 *1 629.595,853.995 sg13_lv_pmos
M$2854 VDD \$25867 \$26450 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2855 r0 *1 620.95,854.02 sg13_lv_pmos
M$2855 VDD \$25867 \$25853 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2856 r0 *1 622.39,854.02 sg13_lv_pmos
M$2856 VDD \$4796 \$26446 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2857 r0 *1 635.87,854.005 sg13_lv_pmos
M$2857 VDD \$26454 \$26920 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2859 r0 *1 637.86,854.02 sg13_lv_pmos
M$2859 VDD \$25840 \$26455 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2860 r0 *1 638.37,854.005 sg13_lv_pmos
M$2860 VDD \$26455 \$26921 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2862 r0 *1 640.39,854.005 sg13_lv_pmos
M$2862 VDD \$26920 \$28308 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2864 r0 *1 617.465,865.11 sg13_lv_pmos
M$2864 VDD \$26953 \$26937 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2866 r0 *1 618.495,865.11 sg13_lv_pmos
M$2866 VDD \$26954 \$26937 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2868 r0 *1 623.525,853.755 sg13_lv_pmos
M$2868 VDD \$25840 \$26447 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2869 r0 *1 624.035,853.755 sg13_lv_pmos
M$2869 VDD \$26446 \$26447 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2870 r0 *1 624.485,854.045 sg13_lv_pmos
M$2870 VDD \$26494 \$26448 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2871 r0 *1 625.535,854.12 sg13_lv_pmos
M$2871 \$26494 \$26446 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2872 r0 *1 626.27,854.12 sg13_lv_pmos
M$2872 VDD \$26448 \$26507 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2873 r0 *1 626.66,854.12 sg13_lv_pmos
M$2873 \$26507 \$26450 \$26494 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2874 r0 *1 627.17,854.12 sg13_lv_pmos
M$2874 \$26494 \$26497 \$26447 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2875 r0 *1 631.725,853.74 sg13_lv_pmos
M$2875 \$26480 \$26497 \$26510 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2876 r0 *1 632.105,853.74 sg13_lv_pmos
M$2876 \$26510 \$26452 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2877 r0 *1 632.715,853.74 sg13_lv_pmos
M$2877 VDD \$26446 \$26452 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2878 r0 *1 633.225,853.74 sg13_lv_pmos
M$2878 VDD \$26480 \$26452 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2879 r0 *1 634.785,853.845 sg13_lv_pmos
M$2879 VDD \$26480 \$26454 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2880 r0 *1 633.765,853.905 sg13_lv_pmos
M$2880 VDD \$26480 \$26453 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2882 r0 *1 631.03,854.03 sg13_lv_pmos
M$2882 \$26448 \$26450 \$26480 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2883 r0 *1 640.7,865.11 sg13_lv_pmos
M$2883 VDD \$26927 \$26938 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2885 r0 *1 641.73,865.11 sg13_lv_pmos
M$2885 VDD \$26926 \$26938 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2887 r0 *1 643.75,865.11 sg13_lv_pmos
M$2887 VDD \$26938 \$26929 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2891 r0 *1 623.374,865.112 sg13_lv_pmos
M$2891 VDD \$26923 \$26924 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2895 r0 *1 626.254,865.112 sg13_lv_pmos
M$2895 VDD \$26924 \$26925 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2899 r0 *1 629.134,865.112 sg13_lv_pmos
M$2899 VDD \$26925 \$26926 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2903 r0 *1 632.714,865.112 sg13_lv_pmos
M$2903 VDD \$26926 \$26142 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2907 r0 *1 636.294,865.112 sg13_lv_pmos
M$2907 VDD \$26142 \$26927 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2911 r0 *1 646.57,865.112 sg13_lv_pmos
M$2911 VDD \$26929 \$26427 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2919 r0 *1 577.495,865.995 sg13_lv_pmos
M$2919 VDD \$26427 \$26956 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2920 r0 *1 578.005,865.995 sg13_lv_pmos
M$2920 VDD \$26920 \$26956 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2921 r0 *1 578.515,865.855 sg13_lv_pmos
M$2921 VDD \$26956 \$26460 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2922 r0 *1 579.805,865.715 sg13_lv_pmos
M$2922 \$26951 \$26920 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2923 r0 *1 580.345,865.855 sg13_lv_pmos
M$2923 VDD \$26427 \$26478 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2924 r0 *1 580.855,865.855 sg13_lv_pmos
M$2924 \$26478 \$26951 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2925 r0 *1 582.565,865.87 sg13_lv_pmos
M$2925 VDD \$25867 \$26426 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2926 r0 *1 599.085,865.995 sg13_lv_pmos
M$2926 VDD \$25867 \$26957 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2927 r0 *1 599.595,865.995 sg13_lv_pmos
M$2927 VDD \$26921 \$26957 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2928 r0 *1 600.105,865.855 sg13_lv_pmos
M$2928 VDD \$26957 \$26461 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2929 r0 *1 601.395,865.715 sg13_lv_pmos
M$2929 \$26952 \$26921 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2930 r0 *1 601.935,865.855 sg13_lv_pmos
M$2930 VDD \$25867 \$26479 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2931 r0 *1 602.445,865.855 sg13_lv_pmos
M$2931 \$26479 \$26952 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2932 r0 *1 604.155,865.87 sg13_lv_pmos
M$2932 VDD \$26427 \$26428 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2933 r0 *1 620.494,870.782 sg13_lv_pmos
M$2933 VDD \$27009 \$26995 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2937 r0 *1 620.494,865.114 sg13_lv_pmos
M$2937 VDD \$26937 \$26923 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2941 r0 *1 623.374,870.782 sg13_lv_pmos
M$2941 VDD \$26995 \$26996 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2945 r0 *1 626.254,870.782 sg13_lv_pmos
M$2945 VDD \$26996 \$26997 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2949 r0 *1 629.134,870.782 sg13_lv_pmos
M$2949 VDD \$26997 \$26998 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2953 r0 *1 632.714,870.782 sg13_lv_pmos
M$2953 VDD \$26998 \$26999 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2957 r0 *1 636.294,870.782 sg13_lv_pmos
M$2957 VDD \$26999 \$26953 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2961 r0 *1 643.505,870.782 sg13_lv_pmos
M$2961 VDD \$27010 \$27001 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2965 r0 *1 613.56,870.787 sg13_lv_pmos
M$2965 VDD \$27008 \$26954 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2967 r0 *1 615.48,870.787 sg13_lv_pmos
M$2967 VDD \$26954 \$26993 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2969 r0 *1 617.465,870.787 sg13_lv_pmos
M$2969 VDD \$26927 \$27009 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2971 r0 *1 618.495,870.787 sg13_lv_pmos
M$2971 VDD \$26993 \$27009 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2973 r0 *1 640.44,870.787 sg13_lv_pmos
M$2973 VDD \$26953 \$27010 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2975 r0 *1 641.47,870.787 sg13_lv_pmos
M$2975 VDD \$26998 \$27010 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2977 r0 *1 646.325,870.788 sg13_lv_pmos
M$2977 VDD \$27001 \$25867 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2985 r0 *1 1056.005,897.48 sg13_lv_pmos
M$2985 \$28306 \$28308 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2986 r0 *1 1056.005,900.99 sg13_lv_pmos
M$2986 \$28334 \$28308 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2987 r0 *1 478.37,933.458 sg13_lv_pmos
M$2987 \$29051 \$29048 \$30346 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $2990 r0 *1 483.435,934.514 sg13_lv_pmos
M$2990 VDD \$29052 \$29048 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2991 r0 *1 438.7,942.5 sg13_lv_pmos
M$2991 VDD \$29422 \$29396 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2993 r0 *1 439.73,942.5 sg13_lv_pmos
M$2993 VDD \$29423 \$29396 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2995 r0 *1 441.615,942.5 sg13_lv_pmos
M$2995 VDD \$29396 \$29397 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2999 r0 *1 444.495,942.5 sg13_lv_pmos
M$2999 VDD \$29397 \$29398 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3003 r0 *1 447.375,942.5 sg13_lv_pmos
M$3003 VDD \$29398 \$29399 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3007 r0 *1 450.255,942.5 sg13_lv_pmos
M$3007 VDD \$29399 \$29400 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3011 r0 *1 453.135,942.5 sg13_lv_pmos
M$3011 VDD \$29400 \$29401 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3015 r0 *1 456.015,942.5 sg13_lv_pmos
M$3015 VDD \$29401 \$29402 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3019 r0 *1 458.97,942.5 sg13_lv_pmos
M$3019 VDD \$29402 \$29403 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3021 r0 *1 460,942.5 sg13_lv_pmos
M$3021 VDD \$29400 \$29403 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3023 r0 *1 461.775,942.5 sg13_lv_pmos
M$3023 VDD \$29403 \$29404 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3027 r0 *1 464.595,942.5 sg13_lv_pmos
M$3027 VDD \$29404 \$29405 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $3035 r0 *1 434.905,948.16 sg13_lv_pmos
M$3035 VDD \$29531 \$29423 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3037 r0 *1 436.825,948.16 sg13_lv_pmos
M$3037 VDD \$29423 \$29492 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3039 r0 *1 438.7,948.16 sg13_lv_pmos
M$3039 VDD \$29492 \$29509 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3041 r0 *1 439.73,948.16 sg13_lv_pmos
M$3041 VDD \$29402 \$29509 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3043 r0 *1 441.615,948.16 sg13_lv_pmos
M$3043 VDD \$29509 \$29494 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3047 r0 *1 444.495,948.16 sg13_lv_pmos
M$3047 VDD \$29494 \$29495 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3051 r0 *1 447.375,948.16 sg13_lv_pmos
M$3051 VDD \$29495 \$29496 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3055 r0 *1 450.255,948.16 sg13_lv_pmos
M$3055 VDD \$29496 \$29497 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3059 r0 *1 453.135,948.16 sg13_lv_pmos
M$3059 VDD \$29497 \$29498 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3063 r0 *1 456.015,948.16 sg13_lv_pmos
M$3063 VDD \$29498 \$29422 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3067 r0 *1 458.97,948.16 sg13_lv_pmos
M$3067 VDD \$29422 \$29510 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3069 r0 *1 460,948.16 sg13_lv_pmos
M$3069 VDD \$29497 \$29510 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3071 r0 *1 461.775,948.16 sg13_lv_pmos
M$3071 VDD \$29510 \$29500 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $3075 r0 *1 464.595,948.16 sg13_lv_pmos
M$3075 VDD \$29500 \$29052 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $3083 r0 *1 477.191,946.747 sg13_lv_pmos
M$3083 \$29485 \$29405 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3084 r0 *1 477.191,945.317 sg13_lv_pmos
M$3084 \$29485 \$29458 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3085 r0 *1 481.99,946.747 sg13_lv_pmos
M$3085 \$29458 \$29485 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3086 r0 *1 481.99,945.317 sg13_lv_pmos
M$3086 \$29458 \$29405 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3087 r0 *1 487.088,945.317 sg13_lv_pmos
M$3087 \$29459 \$29460 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3088 r0 *1 487.088,946.747 sg13_lv_pmos
M$3088 \$29459 \$29458 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3089 r0 *1 492.112,945.305 sg13_lv_pmos
M$3089 \$29460 \$29485 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3090 r0 *1 492.112,946.735 sg13_lv_pmos
M$3090 \$29460 \$29459 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $3091 r0 *1 497.502,945.284 sg13_lv_pmos
M$3091 VDD \$29460 \$29428 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $3092 r0 *1 498.012,945.269 sg13_lv_pmos
M$3092 VDD \$29428 \$29429 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3094 r0 *1 503.36,944.277 sg13_lv_pmos
M$3094 VDD \$4796 \$29392 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3095 r0 *1 504.495,944.012 sg13_lv_pmos
M$3095 VDD \$29460 \$29406 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3096 r0 *1 505.005,944.012 sg13_lv_pmos
M$3096 VDD \$29392 \$29406 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3097 r0 *1 505.455,944.302 sg13_lv_pmos
M$3097 VDD \$29430 \$29407 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $3098 r0 *1 506.505,944.377 sg13_lv_pmos
M$3098 \$29430 \$29392 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3099 r0 *1 507.24,944.377 sg13_lv_pmos
M$3099 VDD \$29407 \$29479 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3100 r0 *1 507.63,944.377 sg13_lv_pmos
M$3100 \$29479 \$29409 \$29430 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3101 r0 *1 508.14,944.377 sg13_lv_pmos
M$3101 \$29430 \$29461 \$29406 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3102 r0 *1 509.84,944.252 sg13_lv_pmos
M$3102 \$29461 \$29409 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3103 r0 *1 510.565,944.252 sg13_lv_pmos
M$3103 VDD \$29052 \$29409 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3104 r0 *1 512.695,943.997 sg13_lv_pmos
M$3104 \$29431 \$29461 \$29481 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3105 r0 *1 513.075,943.997 sg13_lv_pmos
M$3105 \$29481 \$29411 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3106 r0 *1 513.685,943.997 sg13_lv_pmos
M$3106 VDD \$29392 \$29411 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3107 r0 *1 514.195,943.997 sg13_lv_pmos
M$3107 VDD \$29431 \$29411 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $3108 r0 *1 515.755,944.102 sg13_lv_pmos
M$3108 VDD \$29431 \$29413 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $3109 r0 *1 514.735,944.162 sg13_lv_pmos
M$3109 VDD \$29431 \$29412 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3111 r0 *1 512,944.287 sg13_lv_pmos
M$3111 \$29407 \$29409 \$29431 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $3112 r0 *1 516.84,944.262 sg13_lv_pmos
M$3112 VDD \$29413 \$29414 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3114 r0 *1 436.38,963.972 sg13_lv_pmos
M$3114 VDD \$29052 \$30349 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3115 r0 *1 437.455,963.822 sg13_lv_pmos
M$3115 \$30350 \$29414 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $3116 r0 *1 437.995,963.962 sg13_lv_pmos
M$3116 VDD \$29405 \$30351 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3117 r0 *1 438.505,963.962 sg13_lv_pmos
M$3117 \$30351 \$30350 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3118 r0 *1 439.93,964.107 sg13_lv_pmos
M$3118 VDD \$29405 \$30352 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $3119 r0 *1 440.44,964.107 sg13_lv_pmos
M$3119 VDD \$29414 \$30352 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $3120 r0 *1 440.95,963.967 sg13_lv_pmos
M$3120 VDD \$30352 \$30353 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3121 r0 *1 446.163,968.924 sg13_lv_pmos
M$3121 \$30389 \$30349 CORE$12 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $3124 r0 *1 448.83,969.567 sg13_lv_pmos
M$3124 \$30389 \$30351 PAD|VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $3125 r0 *1 454.211,968.657 sg13_lv_pmos
M$3125 \$30340 \$30340 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $3129 r0 *1 458.581,968.642 sg13_lv_pmos
M$3129 \$30343 \$30342 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $3133 r0 *1 465.462,963.972 sg13_lv_pmos
M$3133 VDD \$29405 \$30355 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3134 r0 *1 466.537,963.822 sg13_lv_pmos
M$3134 \$30356 \$29429 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $3135 r0 *1 467.077,963.962 sg13_lv_pmos
M$3135 VDD \$29052 \$30357 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3136 r0 *1 467.587,963.962 sg13_lv_pmos
M$3136 \$30357 \$30356 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3137 r0 *1 469.012,964.107 sg13_lv_pmos
M$3137 VDD \$29052 \$30358 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $3138 r0 *1 469.522,964.107 sg13_lv_pmos
M$3138 VDD \$29429 \$30358 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $3139 r0 *1 470.032,963.967 sg13_lv_pmos
M$3139 VDD \$30358 \$30359 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $3140 r0 *1 475.245,968.924 sg13_lv_pmos
M$3140 \$30390 \$30355 \$30343 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $3143 r0 *1 477.912,969.567 sg13_lv_pmos
M$3143 \$30390 \$30357 PAD|VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $3144 r0 *1 483.293,968.657 sg13_lv_pmos
M$3144 \$30344 \$30344 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $3148 r0 *1 487.663,968.642 sg13_lv_pmos
M$3148 \$30346 \$30345 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $3152 r0 *1 515.9,949.25 sg13_lv_pmos
M$3152 VDD \$29414 \$31708 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $3154 r0 *1 1056.005,997.48 sg13_lv_pmos
M$3154 \$31706 \$31708 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $3155 r0 *1 1056.005,1000.99 sg13_lv_pmos
M$3155 \$31734 \$31708 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $3156 r0 *1 700.255,1056.005 sg13_lv_pmos
M$3156 \$16829 \$32558 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $3157 r0 *1 800.255,1056.005 sg13_lv_pmos
M$3157 \$27008 \$32559 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $3158 r0 *1 900.255,1056.005 sg13_lv_pmos
M$3158 \$29531 \$32560 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $3159 r0 *1 501.765,243.945 sg13_hv_pmos
M$3159 VDD CORE \$4801 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $3160 r0 *1 701.765,243.945 sg13_hv_pmos
M$3160 VDD CORE$1 \$4802 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $3161 r0 *1 801.765,243.945 sg13_hv_pmos
M$3161 VDD CORE$2 \$4803 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $3162 r0 *1 901.765,243.945 sg13_hv_pmos
M$3162 VDD CORE$3 \$4804 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $3163 r0 *1 151.08,285.52 sg13_hv_pmos
M$3163 AVDD \$5435 IN6|PAD AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3203 r0 *1 1141.82,294.58 sg13_hv_pmos
M$3203 IOVDD \$5194 OUT6 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $3219 r0 *1 1068.82,297.64 sg13_hv_pmos
M$3219 \$5742 \$5752 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3220 r0 *1 1068.82,298.47 sg13_hv_pmos
M$3220 IOVDD \$5742 \$5752 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3221 r0 *1 1068.82,299.81 sg13_hv_pmos
M$3221 IOVDD \$5752 \$5927 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3222 r0 *1 1068.82,301.15 sg13_hv_pmos
M$3222 \$5947 \$6134 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3223 r0 *1 1068.82,301.98 sg13_hv_pmos
M$3223 IOVDD \$5947 \$6134 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3224 r0 *1 1068.82,303.32 sg13_hv_pmos
M$3224 IOVDD \$6134 \$5194 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3225 r0 *1 151.08,385.52 sg13_hv_pmos
M$3225 AVDD \$9161 IN5|PAD AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3265 r0 *1 1141.82,394.58 sg13_hv_pmos
M$3265 IOVDD \$9150 OUT5 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $3281 r0 *1 1068.82,397.64 sg13_hv_pmos
M$3281 \$9651 \$9849 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3282 r0 *1 1068.82,398.47 sg13_hv_pmos
M$3282 IOVDD \$9651 \$9849 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3283 r0 *1 1068.82,399.81 sg13_hv_pmos
M$3283 IOVDD \$9849 \$10159 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3284 r0 *1 1068.82,401.15 sg13_hv_pmos
M$3284 \$10175 \$10185 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3285 r0 *1 1068.82,401.98 sg13_hv_pmos
M$3285 IOVDD \$10175 \$10185 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3286 r0 *1 1068.82,403.32 sg13_hv_pmos
M$3286 IOVDD \$10185 \$9150 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3287 r0 *1 151.08,485.52 sg13_hv_pmos
M$3287 AVDD \$13297 IN4|PAD AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3327 r0 *1 1141.82,494.58 sg13_hv_pmos
M$3327 IOVDD \$13286 OUT4 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $3343 r0 *1 1068.82,497.64 sg13_hv_pmos
M$3343 \$13603 \$13787 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3344 r0 *1 1068.82,498.47 sg13_hv_pmos
M$3344 IOVDD \$13603 \$13787 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3345 r0 *1 1068.82,499.81 sg13_hv_pmos
M$3345 IOVDD \$13787 \$13971 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3346 r0 *1 1068.82,501.15 sg13_hv_pmos
M$3346 \$13983 \$13990 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3347 r0 *1 1068.82,501.98 sg13_hv_pmos
M$3347 IOVDD \$13983 \$13990 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3348 r0 *1 1068.82,503.32 sg13_hv_pmos
M$3348 IOVDD \$13990 \$13286 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3349 r0 *1 151.08,585.52 sg13_hv_pmos
M$3349 AVDD \$16712 PAD|VLO AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3389 r0 *1 151.08,685.52 sg13_hv_pmos
M$3389 AVDD \$19878 PAD|VHI AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3429 r0 *1 1125.09,678.44 sg13_hv_pmos
M$3429 IOVDD \$19262 \$19407 IOVDD sg13_hv_pmos W=350.0 L=0.5
* device instance $3479 r0 *1 151.08,785.52 sg13_hv_pmos
M$3479 AVDD \$23953 IN3|PAD AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3519 r0 *1 1141.82,794.58 sg13_hv_pmos
M$3519 IOVDD \$23485 OUT3 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $3535 r0 *1 1068.82,797.64 sg13_hv_pmos
M$3535 \$24420 \$24429 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3536 r0 *1 1068.82,798.47 sg13_hv_pmos
M$3536 IOVDD \$24420 \$24429 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3537 r0 *1 1068.82,799.81 sg13_hv_pmos
M$3537 IOVDD \$24429 \$24435 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3538 r0 *1 1068.82,801.15 sg13_hv_pmos
M$3538 \$24447 \$24454 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3539 r0 *1 1068.82,801.98 sg13_hv_pmos
M$3539 IOVDD \$24447 \$24454 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3540 r0 *1 1068.82,803.32 sg13_hv_pmos
M$3540 IOVDD \$24454 \$23485 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3541 r0 *1 519.105,828.1 sg13_hv_pmos
M$3541 IOVDD \$25328 PAD|VLDO IOVDD sg13_hv_pmos W=1414.0 L=0.44999999999999996
* device instance $3569 r0 *1 497.865,880.705 sg13_hv_pmos
M$3569 IOVDD \$26978 \$26978 IOVDD sg13_hv_pmos W=54.0 L=0.8999999999999999
* device instance $3587 r0 *1 151.08,885.52 sg13_hv_pmos
M$3587 AVDD \$27865 IN2|PAD AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3607 r0 *1 495.265,883.64 sg13_hv_pmos
M$3607 \$26530 \$26530 IOVDD IOVDD sg13_hv_pmos W=1.0 L=5.0
* device instance $3608 r0 *1 497.865,886.92 sg13_hv_pmos
M$3608 IOVDD \$26978 \$26529 IOVDD sg13_hv_pmos W=54.0 L=0.8999999999999999
* device instance $3626 r0 *1 527.575,885.93 sg13_hv_pmos
M$3626 IOVDD \$26919 \$26919 IOVDD sg13_hv_pmos W=36.0 L=0.8999999999999999
* device instance $3632 r0 *1 535.255,885.93 sg13_hv_pmos
M$3632 IOVDD \$26919 \$25328 IOVDD sg13_hv_pmos W=36.0 L=0.8999999999999999
* device instance $3658 r0 *1 1068.82,899.81 sg13_hv_pmos
M$3658 IOVDD \$28320 \$28323 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3659 r0 *1 1068.82,897.64 sg13_hv_pmos
M$3659 \$28307 \$28320 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3660 r0 *1 1068.82,898.47 sg13_hv_pmos
M$3660 IOVDD \$28307 \$28320 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3661 r0 *1 1141.82,894.58 sg13_hv_pmos
M$3661 IOVDD \$27432 OUT2 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $3677 r0 *1 1068.82,901.15 sg13_hv_pmos
M$3677 \$28335 \$28342 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3678 r0 *1 1068.82,901.98 sg13_hv_pmos
M$3678 IOVDD \$28335 \$28342 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3679 r0 *1 1068.82,903.32 sg13_hv_pmos
M$3679 IOVDD \$28342 \$27432 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3680 r0 *1 151.08,985.52 sg13_hv_pmos
M$3680 AVDD \$31321 IN1|PAD AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3720 r0 *1 1141.82,994.58 sg13_hv_pmos
M$3720 IOVDD \$30871 OUT1 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $3736 r0 *1 1068.82,997.64 sg13_hv_pmos
M$3736 \$31707 \$31717 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3737 r0 *1 1068.82,998.47 sg13_hv_pmos
M$3737 IOVDD \$31707 \$31717 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3738 r0 *1 1068.82,999.81 sg13_hv_pmos
M$3738 IOVDD \$31717 \$31723 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3739 r0 *1 1068.82,1001.15 sg13_hv_pmos
M$3739 \$31735 \$31742 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3740 r0 *1 1068.82,1001.98 sg13_hv_pmos
M$3740 IOVDD \$31735 \$31742 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $3741 r0 *1 1068.82,1003.32 sg13_hv_pmos
M$3741 IOVDD \$31742 \$30871 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $3742 r0 *1 701.765,1056.055 sg13_hv_pmos
M$3742 VDD CORE$13 \$32558 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $3743 r0 *1 801.765,1056.055 sg13_hv_pmos
M$3743 VDD CORE$14 \$32559 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $3744 r0 *1 901.765,1056.055 sg13_hv_pmos
M$3744 VDD CORE$15 \$32560 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $3745 r0 *1 278.44,1125.09 sg13_hv_pmos
M$3745 AVDD \$33694 \$33299 AVDD sg13_hv_pmos W=350.0 L=0.5
* device instance $3795 r0 *1 578.44,1125.09 sg13_hv_pmos
M$3795 IOVDD \$33695 \$33300 IOVDD sg13_hv_pmos W=350.0 L=0.5
* device instance $3845 r0 *1 978.44,1125.09 sg13_hv_pmos
M$3845 VDD \$33696 \$33301 VDD sg13_hv_pmos W=350.0 L=0.5
* device instance $3895 r0 *1 385.52,1141.82 sg13_hv_pmos
M$3895 AVDD \$33540 PAD|VREF AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3935 r0 *1 485.52,1148.92 sg13_hv_pmos
M$3935 AVDD \$33541 PAD|VLDO AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3975 r0 *1 264.54,104.19 dantenna
D$3975 VSS VSS dantenna A=35.0028 P=58.08 m=10
* device instance $3979 r0 *1 464.54,104.19 dantenna
D$3979 VSS PAD|RES dantenna A=35.0028 P=58.08 m=2
* device instance $3983 r0 *1 664.54,104.19 dantenna
D$3983 VSS CK4|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $3985 r0 *1 764.54,104.19 dantenna
D$3985 VSS CK5|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $3987 r0 *1 864.54,104.19 dantenna
D$3987 VSS CK6|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $3991 r0 *1 100.44,400 dantenna
D$3991 VSS IN5|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $3992 r0 *1 100.44,300 dantenna
D$3992 VSS IN6|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $3995 r0 *1 222.54,417.63 dantenna
D$3995 VSS CORE$5 dantenna A=1.984 P=7.48 m=1
* device instance $3996 r0 *1 222.54,317.63 dantenna
D$3996 VSS CORE$4 dantenna A=1.984 P=7.48 m=1
* device instance $3997 r0 *1 505.225,222.54 dantenna
D$3997 VSS CORE dantenna A=1.984 P=7.48 m=1
* device instance $3998 r0 *1 705.225,222.54 dantenna
D$3998 VSS CORE$1 dantenna A=1.984 P=7.48 m=1
* device instance $3999 r0 *1 805.225,222.54 dantenna
D$3999 VSS CORE$2 dantenna A=1.984 P=7.48 m=1
* device instance $4000 r0 *1 905.225,222.54 dantenna
D$4000 VSS CORE$3 dantenna A=1.984 P=7.48 m=1
* device instance $4001 r0 *1 1195.06,300 dantenna
D$4001 VSS OUT6 dantenna A=35.0028 P=58.08 m=2
* device instance $4002 r0 *1 1195.06,400 dantenna
D$4002 VSS OUT5 dantenna A=35.0028 P=58.08 m=2
* device instance $4005 r0 *1 1207.17,377.975 dantenna
D$4005 VSS \$10159 dantenna A=0.192 P=1.88 m=1
* device instance $4006 r0 *1 1207.17,277.975 dantenna
D$4006 VSS \$5927 dantenna A=0.192 P=1.88 m=1
* device instance $4007 r0 *1 1207.17,477.975 dantenna
D$4007 VSS \$13971 dantenna A=0.192 P=1.88 m=1
* device instance $4008 r0 *1 100.44,500 dantenna
D$4008 VSS IN4|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $4010 r0 *1 1195.06,500 dantenna
D$4010 VSS OUT4 dantenna A=35.0028 P=58.08 m=2
* device instance $4012 r0 *1 222.54,517.63 dantenna
D$4012 VSS CORE$6 dantenna A=1.984 P=7.48 m=1
* device instance $4015 r0 *1 100.44,600 dantenna
D$4015 VSS PAD|VLO dantenna A=35.0028 P=58.08 m=2
* device instance $4017 r0 *1 222.54,617.63 dantenna
D$4017 VSS CORE$7 dantenna A=1.984 P=7.48 m=1
* device instance $4018 r0 *1 1192.65,664.765 dantenna
D$4018 VSS \$19407 dantenna A=0.192 P=1.88 m=1
* device instance $4019 r0 *1 100.44,700 dantenna
D$4019 VSS PAD|VHI dantenna A=35.0028 P=58.08 m=2
* device instance $4021 r0 *1 222.54,717.63 dantenna
D$4021 VSS CORE$8 dantenna A=1.984 P=7.48 m=1
* device instance $4022 r0 *1 1207.17,777.975 dantenna
D$4022 VSS \$24435 dantenna A=0.192 P=1.88 m=1
* device instance $4023 r0 *1 100.44,800 dantenna
D$4023 VSS IN3|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $4025 r0 *1 1195.06,800 dantenna
D$4025 VSS OUT3 dantenna A=35.0028 P=58.08 m=2
* device instance $4027 r0 *1 222.54,817.63 dantenna
D$4027 VSS CORE$9 dantenna A=1.984 P=7.48 m=1
* device instance $4028 r0 *1 1207.17,877.975 dantenna
D$4028 VSS \$28323 dantenna A=0.192 P=1.88 m=1
* device instance $4029 r0 *1 100.44,900 dantenna
D$4029 VSS IN2|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $4031 r0 *1 1195.06,900 dantenna
D$4031 VSS OUT2 dantenna A=35.0028 P=58.08 m=2
* device instance $4033 r0 *1 222.54,917.63 dantenna
D$4033 VSS CORE$11 dantenna A=1.984 P=7.48 m=1
* device instance $4034 r0 *1 1207.17,977.975 dantenna
D$4034 VSS \$31723 dantenna A=0.192 P=1.88 m=1
* device instance $4035 r0 *1 100.44,1000 dantenna
D$4035 VSS IN1|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $4037 r0 *1 1195.06,1000 dantenna
D$4037 VSS OUT1 dantenna A=35.0028 P=58.08 m=2
* device instance $4039 r0 *1 222.54,1017.63 dantenna
D$4039 VSS CORE$12 dantenna A=1.984 P=7.48 m=1
* device instance $4040 r0 *1 417.63,1077.46 dantenna
D$4040 VSS CORE$10 dantenna A=1.984 P=7.48 m=1
* device instance $4041 r0 *1 517.63,1077.46 dantenna
D$4041 VSS CORE$16 dantenna A=1.984 P=7.48 m=1
* device instance $4042 r0 *1 705.225,1077.46 dantenna
D$4042 VSS CORE$13 dantenna A=1.984 P=7.48 m=1
* device instance $4043 r0 *1 805.225,1077.46 dantenna
D$4043 VSS CORE$14 dantenna A=1.984 P=7.48 m=1
* device instance $4044 r0 *1 905.225,1077.46 dantenna
D$4044 VSS CORE$15 dantenna A=1.984 P=7.48 m=1
* device instance $4045 r0 *1 664.54,1195.81 dantenna
D$4045 VSS CK3|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $4047 r0 *1 764.54,1195.81 dantenna
D$4047 VSS CK2|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $4049 r0 *1 864.54,1195.81 dantenna
D$4049 VSS CK1|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $4051 r0 *1 264.765,1192.65 dantenna
D$4051 VSS \$33299 dantenna A=0.192 P=1.88 m=1
* device instance $4052 r0 *1 400,1195.06 dantenna
D$4052 VSS PAD|VREF dantenna A=35.0028 P=58.08 m=2
* device instance $4053 r0 *1 500,1195.06 dantenna
D$4053 VSS PAD|VLDO dantenna A=35.0028 P=58.08 m=2
* device instance $4054 r0 *1 564.765,1192.65 dantenna
D$4054 VSS \$33300 dantenna A=0.192 P=1.88 m=1
* device instance $4055 r0 *1 964.765,1192.65 dantenna
D$4055 VSS \$33301 dantenna A=0.192 P=1.88 m=1
* device instance $4058 r0 *1 264.54,163.19 dpantenna
D$4058 VSS AVDD dpantenna A=35.0028 P=58.08 m=4
* device instance $4062 r0 *1 464.54,163.19 dpantenna
D$4062 PAD|RES IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4064 r0 *1 564.54,163.19 dpantenna
D$4064 VSS IOVDD dpantenna A=35.0028 P=58.08 m=6
* device instance $4066 r0 *1 664.54,163.19 dpantenna
D$4066 CK4|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4068 r0 *1 764.54,163.19 dpantenna
D$4068 CK5|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4070 r0 *1 864.54,163.19 dpantenna
D$4070 CK6|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4074 r0 *1 227.51,315.46 dpantenna
D$4074 CORE$4 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4075 r0 *1 227.51,415.46 dpantenna
D$4075 CORE$5 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4076 r0 *1 227.51,515.46 dpantenna
D$4076 CORE$6 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4077 r0 *1 227.51,615.46 dpantenna
D$4077 CORE$7 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4078 r0 *1 227.51,715.46 dpantenna
D$4078 CORE$8 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4079 r0 *1 227.51,815.46 dpantenna
D$4079 CORE$9 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4080 r0 *1 227.51,915.46 dpantenna
D$4080 CORE$11 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4081 r0 *1 227.51,1015.46 dpantenna
D$4081 CORE$12 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4082 r0 *1 415.46,1072.49 dpantenna
D$4082 CORE$10 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4083 r0 *1 515.46,1072.49 dpantenna
D$4083 CORE$16 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4084 r0 *1 503.055,227.51 dpantenna
D$4084 CORE IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4085 r0 *1 703.055,227.51 dpantenna
D$4085 CORE$1 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4086 r0 *1 803.055,227.51 dpantenna
D$4086 CORE$2 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4087 r0 *1 903.055,227.51 dpantenna
D$4087 CORE$3 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4088 r0 *1 703.055,1072.49 dpantenna
D$4088 CORE$13 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4089 r0 *1 803.055,1072.49 dpantenna
D$4089 CORE$14 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4090 r0 *1 903.055,1072.49 dpantenna
D$4090 CORE$15 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $4091 r0 *1 1138.81,277.975 dpantenna
D$4091 \$5194 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $4092 r0 *1 135.96,300 dpantenna
D$4092 IN6|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4094 r0 *1 1159.54,300 dpantenna
D$4094 OUT6 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4096 r0 *1 135.96,400 dpantenna
D$4096 IN5|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4098 r0 *1 1138.81,377.975 dpantenna
D$4098 \$9150 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $4099 r0 *1 1159.54,400 dpantenna
D$4099 OUT5 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4101 r0 *1 135.96,500 dpantenna
D$4101 IN4|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4103 r0 *1 1138.81,477.975 dpantenna
D$4103 \$13286 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $4104 r0 *1 1159.54,500 dpantenna
D$4104 OUT4 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4106 r0 *1 135.96,600 dpantenna
D$4106 PAD|VLO AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4110 r0 *1 135.96,700 dpantenna
D$4110 PAD|VHI AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4112 r0 *1 1138.81,777.975 dpantenna
D$4112 \$23485 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $4113 r0 *1 135.96,800 dpantenna
D$4113 IN3|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4115 r0 *1 1159.54,800 dpantenna
D$4115 OUT3 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4117 r0 *1 135.96,900 dpantenna
D$4117 IN2|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4119 r0 *1 1138.81,877.975 dpantenna
D$4119 \$27432 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $4120 r0 *1 1159.54,900 dpantenna
D$4120 OUT2 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4122 r0 *1 135.96,1000 dpantenna
D$4122 IN1|PAD AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4124 r0 *1 1138.81,977.975 dpantenna
D$4124 \$30871 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $4125 r0 *1 1159.54,1000 dpantenna
D$4125 OUT1 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4127 r0 *1 664.54,1136.81 dpantenna
D$4127 CK3|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4129 r0 *1 764.54,1136.81 dpantenna
D$4129 CK2|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4131 r0 *1 864.54,1136.81 dpantenna
D$4131 CK1|PAD IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4133 r0 *1 400,1159.54 dpantenna
D$4133 PAD|VREF AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4135 r0 *1 500,1159.54 dpantenna
D$4135 PAD|VLDO AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $4137 r0 *1 500.685,221.11 rppd
R$4137 PAD|RES CORE rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4138 r0 *1 700.685,221.11 rppd
R$4138 CK4|PAD CORE$1 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4139 r0 *1 800.685,221.11 rppd
R$4139 CK5|PAD CORE$2 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4140 r0 *1 900.685,221.11 rppd
R$4140 CK6|PAD CORE$3 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4141 r0 *1 88.75,326.305 rppd
R$4141 VSS \$5434 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4142 r0 *1 147.75,326.305 rppd
R$4142 AVDD \$5435 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4143 r0 *1 221.11,313.09 rppd
R$4143 IN6|PAD CORE$4 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4144 r0 *1 88.75,426.305 rppd
R$4144 VSS \$9160 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4145 r0 *1 147.75,426.305 rppd
R$4145 AVDD \$9161 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4146 r0 *1 221.11,413.09 rppd
R$4146 IN5|PAD CORE$5 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4147 r0 *1 88.75,526.305 rppd
R$4147 VSS \$13296 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4148 r0 *1 147.75,526.305 rppd
R$4148 AVDD \$13297 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4149 r0 *1 221.11,513.09 rppd
R$4149 IN4|PAD CORE$6 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4150 r0 *1 88.75,626.305 rppd
R$4150 VSS \$16711 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4151 r0 *1 147.75,626.305 rppd
R$4151 AVDD \$16712 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4152 r0 *1 221.11,613.09 rppd
R$4152 PAD|VLO CORE$7 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4153 r0 *1 1161.29,678.875 rppd
R$4153 IOVDD \$19262 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $4154 r0 *1 221.11,713.09 rppd
R$4154 PAD|VHI CORE$8 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4155 r0 *1 88.75,726.305 rppd
R$4155 VSS \$19877 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4156 r0 *1 147.75,726.305 rppd
R$4156 AVDD \$19878 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4157 r0 *1 88.75,826.305 rppd
R$4157 VSS \$23952 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4158 r0 *1 147.75,826.305 rppd
R$4158 AVDD \$23953 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4159 r0 *1 221.11,813.09 rppd
R$4159 IN3|PAD CORE$9 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4160 r0 *1 221.11,913.09 rppd
R$4160 IN2|PAD CORE$11 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4161 r0 *1 88.75,926.305 rppd
R$4161 VSS \$27864 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4162 r0 *1 147.75,926.305 rppd
R$4162 AVDD \$27865 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4163 r0 *1 88.75,1026.305 rppd
R$4163 VSS \$31320 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4164 r0 *1 147.75,1026.305 rppd
R$4164 AVDD \$31321 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4165 r0 *1 221.11,1013.09 rppd
R$4165 IN1|PAD CORE$12 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4166 r0 *1 413.09,1076.03 rppd
R$4166 CORE$10 PAD|VREF rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4167 r0 *1 513.09,1076.03 rppd
R$4167 CORE$16 PAD|VLDO rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4168 r0 *1 700.685,1076.03 rppd
R$4168 CORE$13 CK3|PAD rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4169 r0 *1 800.685,1076.03 rppd
R$4169 CORE$14 CK2|PAD rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4170 r0 *1 900.685,1076.03 rppd
R$4170 CORE$15 CK1|PAD rppd w=1 l=2 ps=0 b=0 m=1
* device instance $4171 r0 *1 278.875,1161.29 rppd
R$4171 AVDD \$33694 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $4172 r0 *1 426.305,1138.49 rppd
R$4172 \$33540 AVDD rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4173 r0 *1 526.305,1138.49 rppd
R$4173 \$33541 AVDD rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $4174 r0 *1 578.875,1161.29 rppd
R$4174 IOVDD \$33695 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $4175 r0 *1 978.875,1161.29 rppd
R$4175 VDD \$33696 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $4176 r0 *1 426.305,1206.85 rppd
R$4176 \$34430 VSS rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4177 r0 *1 526.305,1206.85 rppd
R$4177 \$34431 VSS rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $4178 r0 *1 506.575,859.565 rhigh
R$4178 VSS \$26955 rhigh w=0.5 l=0.96 ps=0 b=0 m=2
* device instance $4182 r0 *1 543.535,883.575 rhigh
R$4182 \$25328 \$25329 rhigh w=0.5 l=3.84 ps=0 b=0 m=1
* device instance $4184 r0 *1 463.265,300.165 cap_cmim
C$4184 \$6118 \$6133 cap_cmim w=8.16 l=8.16 m=1
* device instance $4185 r0 *1 463.27,309.855 cap_cmim
C$4185 \$6145 \$6117 cap_cmim w=8.16 l=8.16 m=1
* device instance $4186 r0 *1 455.04,311.655 cap_cmim
C$4186 \$6133 \$6193 cap_cmim w=5.77 l=5.77 m=1
* device instance $4187 r0 *1 438.16,318.59 cap_cmim
C$4187 \$6783 \$6774 cap_cmim w=8.16 l=8.16 m=1
* device instance $4188 r0 *1 438.165,328.28 cap_cmim
C$4188 \$7040 \$6197 cap_cmim w=8.16 l=8.16 m=1
* device instance $4189 r0 *1 429.935,330.08 cap_cmim
C$4189 \$6774 \$7314 cap_cmim w=5.77 l=5.77 m=1
* device instance $4190 r0 *1 439.894,391.265 cap_cmim
C$4190 \$9622 \$9623 cap_cmim w=8.16 l=8.16 m=1
* device instance $4191 r0 *1 449.03,330.495 cap_cmim
C$4191 \$7364 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $4192 r0 *1 492.368,391.265 cap_cmim
C$4192 \$9625 \$9624 cap_cmim w=8.16 l=8.16 m=1
* device instance $4193 r0 *1 449.469,391.27 cap_cmim
C$4193 \$9623 \$9634 cap_cmim w=5.77 l=5.77 m=1
* device instance $4194 r0 *1 457.713,410.953 cap_cmim
C$4194 \$10369 \$10410 cap_cmim w=8.16 l=8.16 m=1
* device instance $4195 r0 *1 474.549,410.953 cap_cmim
C$4195 \$10370 \$10411 cap_cmim w=8.16 l=8.16 m=1
* device instance $4196 r0 *1 485.183,391.27 cap_cmim
C$4196 \$9624 \$9848 cap_cmim w=5.77 l=5.77 m=1
* device instance $4197 r0 *1 471.467,445.302 cap_cmim
C$4197 \$11659 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $4198 r0 *1 473.164,512.175 cap_cmim
C$4198 \$14122 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $4199 r0 *1 430.955,540.411 cap_cmim
C$4199 \$15333 \$15336 cap_cmim w=5.77 l=5.77 m=1
* device instance $4200 r0 *1 465.955,540.411 cap_cmim
C$4200 \$15334 \$15076 cap_cmim w=5.77 l=5.77 m=1
* device instance $4201 r0 *1 439.56,542.231 cap_cmim
C$4201 \$15047 \$15333 cap_cmim w=8.16 l=8.16 m=1
* device instance $4202 r0 *1 474.56,542.231 cap_cmim
C$4202 \$15049 \$15334 cap_cmim w=8.16 l=8.16 m=1
* device instance $4203 r0 *1 443.88,615.55 cap_cmim
C$4203 \$17393 \$17495 cap_cmim w=5.77 l=5.77 m=1
* device instance $4204 r0 *1 450.88,542.236 cap_cmim
C$4204 \$15048 \$15341 cap_cmim w=8.16 l=8.16 m=1
* device instance $4205 r0 *1 479.935,615.55 cap_cmim
C$4205 \$17394 \$17540 cap_cmim w=5.77 l=5.77 m=1
* device instance $4206 r0 *1 485.88,542.236 cap_cmim
C$4206 \$14121 \$15335 cap_cmim w=8.16 l=8.16 m=1
* device instance $4207 r0 *1 509.38,615.465 cap_cmim
C$4207 \$17662 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $4208 r0 *1 430.19,624.19 cap_cmim
C$4208 \$17673 \$17496 cap_cmim w=8.16 l=8.16 m=1
* device instance $4209 r0 *1 466.245,624.19 cap_cmim
C$4209 \$17674 \$17497 cap_cmim w=8.16 l=8.16 m=1
* device instance $4210 r0 *1 441.11,625.165 cap_cmim
C$4210 \$17412 \$17393 cap_cmim w=8.16 l=8.16 m=1
* device instance $4211 r0 *1 477.165,625.165 cap_cmim
C$4211 \$17413 \$17394 cap_cmim w=8.16 l=8.16 m=1
* device instance $4212 r0 *1 429.41,826.865 cap_cmim
C$4212 \$25329 PAD|VLDO cap_cmim w=60 l=60 m=1
* device instance $4213 r0 *1 429.41,682.847 cap_cmim
C$4213 VSS PAD|VLDO cap_cmim w=140 l=225 m=1
* device instance $4214 r0 *1 623.755,834.77 cap_cmim
C$4214 \$25487 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $4215 r0 *1 576.305,835.415 cap_cmim
C$4215 \$25489 \$25851 cap_cmim w=8.16 l=8.16 m=1
* device instance $4216 r0 *1 587.54,835.275 cap_cmim
C$4216 \$25485 \$25833 cap_cmim w=8.16 l=8.16 m=1
* device instance $4217 r0 *1 597.895,835.415 cap_cmim
C$4217 \$25490 \$25852 cap_cmim w=8.16 l=8.16 m=1
* device instance $4218 r0 *1 609.13,835.275 cap_cmim
C$4218 \$25486 \$25822 cap_cmim w=8.16 l=8.16 m=1
* device instance $4219 r0 *1 576.185,848.635 cap_cmim
C$4219 \$25851 \$25848 cap_cmim w=5.77 l=5.77 m=1
* device instance $4220 r0 *1 597.775,848.635 cap_cmim
C$4220 \$25852 \$25849 cap_cmim w=5.77 l=5.77 m=1
* device instance $4221 r0 *1 484.503,930.308 cap_cmim
C$4221 \$29051 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $4222 r0 *1 435.608,966.963 cap_cmim
C$4222 \$30354 \$30389 cap_cmim w=5.77 l=5.77 m=1
* device instance $4223 r0 *1 464.69,966.963 cap_cmim
C$4223 \$30360 \$30390 cap_cmim w=5.77 l=5.77 m=1
* device instance $4224 r0 *1 434.36,974.656 cap_cmim
C$4224 \$30342 \$30354 cap_cmim w=8.16 l=8.16 m=1
* device instance $4225 r0 *1 463.442,974.656 cap_cmim
C$4225 \$30345 \$30360 cap_cmim w=8.16 l=8.16 m=1
* device instance $4226 r0 *1 450.71,975.898 cap_cmim
C$4226 \$30341 \$30343 cap_cmim w=8.16 l=8.16 m=1
* device instance $4227 r0 *1 479.792,975.898 cap_cmim
C$4227 \$30361 \$30346 cap_cmim w=8.16 l=8.16 m=1
.ENDS UHEE628_S2024

* Extracted by KLayout with SG13G2 LVS runset on : 29/04/2024 22:26

* cell sg13g2_SecondaryProtection
* pin CORE
* pin PAD
* pin IOVDD
* pin IOVSS
.SUBCKT sg13g2_SecondaryProtection CORE PAD IOVDD IOVSS
* device instance $1 r0 *1 5.48,2.37 dantenna
D$1 IOVSS CORE dantenna A=1.984 P=7.48 m=1
* device instance $2 r0 *1 3.31,7.34 dpantenna
D$2 CORE IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3 r0 *1 0.94,0.94 res_rppd
R$3 PAD CORE res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0 ps=0.0
+ m=1.0
.ENDS sg13g2_SecondaryProtection

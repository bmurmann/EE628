* Extracted by KLayout with SG13G2 LVS runset on : 03/05/2024 02:13

* cell sg13g2_LevelDown
.SUBCKT sg13g2_LevelDown
* net 1 CORE
* net 2 sub!
* net 3 sub!
* net 4 PAD
* net 5 IOVSS
* net 6 rppd r=793.834
* net 7 dant
* net 12 IOVDD
* net 13 dpant
* net 25 sub!
* device instance $1 r0 *1 0.51,10.505 sg13_lv_nmos
M$1 17 18 25 25 sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $2 r0 *1 2.02,10.555 sg13_hv_nmos
M$2 25 1 18 25 sg13_hv_nmos W=2.6499999999999995 L=0.4499999999999999
* device instance $3 r0 *1 0.51,15.495 sg13_lv_pmos
M$3 17 18 21 21 sg13_lv_pmos W=4.749999999999999 L=0.12999999999999998
* device instance $4 r0 *1 2.02,15.445 sg13_hv_pmos
M$4 21 1 18 21 sg13_hv_pmos W=4.6499999999999995 L=0.44999999999999984
* device instance $5 r0 *1 5.48,-5.96 dantenna
D$5 25 1 dantenna A=1.984 P=7.48 m=1
* device instance $6 r0 *1 3.31,-0.99 dpantenna
D$6 1 9 dpantenna A=3.1872 P=11.24 m=1
* device instance $7 r0 *1 0.94,-7.39 rppd
R$7 4 1 rppd w=1 l=2 ps=0 b=0 m=1
.ENDS sg13g2_LevelDown

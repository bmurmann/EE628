** sch_path: /foss/designs/EE628_template/Team_2.sch
.subckt Team_2 vlo vhi vdda vssa iovdd vref vin dd res clkin
*.PININFO clkin:I res:I dd:O vlo:I vssa:I vhi:I vin:I iovdd:I vref:I vdda:B
x1 vmid res p1e p1 p2 vhi vdda vin vssa dd vlo vout1 Stage_T2
x3 p1e clkin p1 p2 p2e ClockGen_T2
x4 vdda p2 net1 dd vmid res vssa p1 vout2 comparator_latch_T2
M2 vmid vmid vdda vdda sg13_lv_pmos L=1.5u W=10u ng=4 m=1
M5 vmid vmid vssa vssa sg13_lv_nmos L=1.5u W=2.5u ng=1 m=1
x5 iovdd vref vdda vssa Team2_LDO_updt
x2 vmid res p2e p2 p1 vhi vdda vout1 vssa net1 vlo vout2 Stage_T2
.ends

* expanding   symbol:  /foss/designs/EE_628_final/Stage_T2.sym # of pins=12
** sym_path: /foss/designs/EE_628_final/Stage_T2.sym
** sch_path: /foss/designs/EE_628_final/Stage_T2.sch
.subckt Stage_T2 vmid res pse ps pr vhi vdda vin vssa d vlo vout
*.PININFO vin:I ps:I pse:I vout:O vmid:B res:I pr:I vdda:B vssa:B vhi:B d:I vlo:B
M3 vout vx3 vdda vdda sg13_lv_pmos L=1.5u W=10u ng=4 m=1
M4 vout vx3 vssa vssa sg13_lv_nmos L=1.5u W=2.5u ng=1 m=1
M1 vx4 pr vx2 vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M6 vx4 ps vx3 vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M7 vx2 pse vmid vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M8 vout res vx4 vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M9 vx1 gn vlo vssa sg13_lv_nmos L=.13u W=0.5u ng=1 m=1
M10 vx1 ps vin vssa sg13_lv_nmos L=0.13u W=2u ng=3 m=1
M11 vx1 psb vin vdda sg13_lv_pmos L=0.13u W=6u ng=1 m=1
x3 ps VDD VSS psb sg13g2_inv_1
M2 vx1 gp vhi vdda sg13_lv_pmos L=0.13u W=1.5u ng=1 m=1
x1 d pr VDD VSS gp sg13g2_nand2b_1
x2 pr d VDD VSS gn sg13g2_and2_1
XC1 vx2 vx1 cap_cmim W=5.77e-6 L=5.77e-6 MF=1
XC2 vx4 vout cap_cmim W=8.16e-6 L=8.16e-6 MF=1
XC3 vx3 vx2 cap_cmim W=8.16e-6 L=8.16e-6 MF=1
.ends


* expanding   symbol:  /foss/designs/EE628_template/ClockGen_T2.sym # of pins=5
** sym_path: /foss/designs/EE628_template/ClockGen_T2.sym
** sch_path: /foss/designs/EE628_template/ClockGen_T2.sch
.subckt ClockGen_T2 p1e clkIn p1 p2 p2e
*.PININFO clkIn:I p1:O p1e:O p2:O p2e:O
x3 net1 net3 VDD VSS net13 sg13g2_nand2_2
x4 net2 net4 VDD VSS net5 sg13g2_nand2_2
x17 net14 net3 VDD VSS net15 sg13g2_nand2_2
x18 net12 net4 VDD VSS net17 sg13g2_nand2_2
x6 net10 VDD VSS net11 sg13g2_inv_4
x7 net11 VDD VSS net12 sg13g2_inv_4
x8 net12 VDD VSS p1e sg13g2_inv_4
x11 net7 VDD VSS net8 sg13g2_inv_4
x12 net8 VDD VSS net14 sg13g2_inv_4
x13 net14 VDD VSS p2e sg13g2_inv_4
x14 p2e VDD VSS net3 sg13g2_inv_4
x15 p1e VDD VSS net4 sg13g2_inv_4
x16 net17 VDD VSS net18 sg13g2_inv_4
x19 net15 VDD VSS net16 sg13g2_inv_4
x20 net18 VDD VSS p1 sg13g2_inv_8
x21 net16 VDD VSS p2 sg13g2_inv_8
x1 net2 VDD VSS net1 sg13g2_inv_2
x2 clkIn VDD VSS net2 sg13g2_inv_2
x5 net5 VDD VSS net6 sg13g2_inv_4
x9 net6 VDD VSS net7 sg13g2_inv_4
x10 net13 VDD VSS net9 sg13g2_inv_4
x23 net9 VDD VSS net10 sg13g2_inv_4
.ends


* expanding   symbol:  /foss/designs/EE_628_final/comparator_latch_T2.sym # of pins=9
** sym_path: /foss/designs/EE_628_final/comparator_latch_T2.sym
** sch_path: /foss/designs/EE_628_final/comparator_latch_T2.sch
.subckt comparator_latch_T2 vdda pc d dd vinp res vssa ps vinm
*.PININFO vdda:B vssa:B pc:I vinp:I vinm:I ps:I dd:O d:O res:I
M1 d2p pc d1p vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M3 out1m pc vdda vdda sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M4 out1m out1p vdda vdda sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M5 out1m out1p d2p vssa sg13_lv_nmos L=0.13u W=2.0u ng=1 m=1
M6 d1p vinp vssa vssa sg13_lv_nmos L=1u W=2.0u ng=1 m=1
M2 out1p out1m vdda vdda sg13_lv_pmos L=0.13u W=4.0u ng=1 m=1
M7 out1p pc vdda vdda sg13_lv_pmos L=0.13u W=4.0u ng=1 m=1
M8 d2m pc d1m vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M9 out1p out1m d2m vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M10 d1m vinm_samp vssa vssa sg13_lv_nmos L=1u W=2.0u ng=1 m=1
M11 d2p2 out1p VSS VSS sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M12 net1 out1p VDD VDD sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M13 net1 net2 VDD VDD sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M14 net1 net2 d2p2 VSS sg13_lv_nmos L=0.13u W=2.0u ng=1 m=1
M16 net2 net1 VDD VDD sg13_lv_pmos L=0.13u W=4.0u ng=1 m=1
M17 net2 out1m VDD VDD sg13_lv_pmos L=0.13u W=4.0u ng=1 m=1
M18 d2m2 out1m VSS VSS sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M19 net2 net1 d2m2 VSS sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M15 vinm_samp ps vinm vssa sg13_lv_nmos L=0.13u W=2.0u ng=1 m=1
M20 vinm_samp net3 vinm vdda sg13_lv_pmos L=0.13u W=4u ng=1 m=1
x1 ps VDD VSS net3 sg13g2_inv_1
x2 net2 VDD VSS d sg13g2_buf_2
x3 ps net2 net5 net6 net4 VDD VSS sg13g2_dfrbp_2
x4 res VDD VSS net4 sg13g2_inv_1
XC1 vinm_samp vssa cap_cmim W=5.77e-6 L=5.77e-6 MF=1
x5 net5 VDD VSS dd sg13g2_inv_1
.ends


* expanding   symbol:  /foss/designs/EE_628_final/Team2_LDO_updt.sym # of pins=4
** sym_path: /foss/designs/EE_628_final/Team2_LDO_updt.sym
** sch_path: /foss/designs/EE_628_final/Team2_LDO_updt.sch
.subckt Team2_LDO_updt Vin Vref Vout VSS
*.PININFO Vin:I Vref:I Vout:O VSS:I
XC3 Vout VSS cap_cmim W=140.0e-6 L=225.0e-6 MF=1
M1 Vout Verr Vin Vin sg13_hv_pmos L=0.45u W=1.414m ng=1 m=1
XC4 Vout net1 cap_cmim W=60.0e-6 L=60.0e-6 MF=1
x1 Vin Verr Vout Vref VSS Team2_DiffAmp_Ref
XR4 Verr net1 rhigh w=0.5e-6 l=5*0.96e-6 m=1 b=0
.ends


* expanding   symbol:  /foss/designs/EE_628_final/Team2_DiffAmp_Ref.sym # of pins=5
** sym_path: /foss/designs/EE_628_final/Team2_DiffAmp_Ref.sym
** sch_path: /foss/designs/EE_628_final/Team2_DiffAmp_Ref.sch
.subckt Team2_DiffAmp_Ref VDD Vout Vp Vm VSS
*.PININFO Vout:O Vm:I Vp:I VDD:I VSS:I
M6 vstart vstart VDD VDD sg13_hv_pmos L=5u W=1.0u ng=1 m=1
M1 vbp vstart VSS VSS sg13_hv_nmos L=0.45u W=1.0u ng=1 m=1
M9 vstart vbn VSS VSS sg13_hv_nmos L=0.9u W=33u ng=1 m=1
M4 vbp vbn net1 VSS sg13_hv_nmos L=0.9u W=178u ng=1 m=1
M13 vbn vbn VSS VSS sg13_hv_nmos L=0.9u W=33u ng=1 m=1
M5 vbp vbp VDD VDD sg13_hv_pmos L=0.9u W=54u ng=1 m=1
M10 vbn vbp VDD VDD sg13_hv_pmos L=0.9u W=54u ng=1 m=1
XR4 VSS net1 rhigh w=0.5e-6 l=0.96e-6 m=2 b=0
M14 Vout net2 VDD VDD sg13_hv_pmos L=0.9u W=36u ng=1 m=1
M16 net2 net2 VDD VDD sg13_hv_pmos L=0.9u W=36u ng=1 m=1
M17 net2 Vp net3 VSS sg13_hv_nmos L=0.9u W=136.5u ng=1 m=1
M18 Vout Vm net3 VSS sg13_hv_nmos L=0.9u W=136.5u ng=1 m=1
M19 net3 vbn VSS VSS sg13_hv_nmos L=0.9u W=33u ng=1 m=1
.ends

.GLOBAL VDD
.GLOBAL VSS
.end

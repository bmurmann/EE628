* Extracted by KLayout with SG13G2 LVS runset on : 02/05/2024 06:31

* cell sg13g2_RCClampResistor
.SUBCKT sg13g2_RCClampResistor
* net 15 rpnd r=5238.986
* net 16 rpnd r=5238.986
* net 17 rpnd r=5238.986
* net 18 rpnd r=5238.986
* net 19 rpnd r=5238.986
* net 20 rpnd r=5238.986
* net 21 rpnd r=5238.986
* net 22 rpnd r=5238.986
* net 23 rpnd r=5238.986
* net 24 rpnd r=5238.986
* net 25 rpnd r=5238.986
* net 26 rpnd r=5238.986
* net 27 rpnd r=5238.986
* net 28 rpnd r=5238.986
* net 29 rpnd r=5238.986
* net 30 rpnd r=5238.986
* net 31 rpnd r=5238.986
* net 32 rpnd r=5238.986
* net 33 rpnd r=5238.986
* net 34 rpnd r=5238.986
* net 35 rpnd r=5238.986
* net 36 rpnd r=5238.986
* net 37 rpnd r=5238.986
* net 38 rpnd r=5238.986
* net 39 rpnd r=5238.986
* net 40 rpnd r=5238.986
* net 54 sub!
* device instance $1 r0 *1 0,0 res_rppd
R$1 1 41 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $2 r0 *1 1.65,0 res_rppd
R$2 2 41 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $3 r0 *1 3.3,0 res_rppd
R$3 2 42 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $4 r0 *1 4.95,0 res_rppd
R$4 3 42 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $5 r0 *1 6.6,0 res_rppd
R$5 3 43 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $6 r0 *1 8.25,0 res_rppd
R$6 4 43 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $7 r0 *1 9.9,0 res_rppd
R$7 4 44 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $8 r0 *1 11.55,0 res_rppd
R$8 5 44 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $9 r0 *1 13.2,0 res_rppd
R$9 5 45 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $10 r0 *1 14.85,0 res_rppd
R$10 6 45 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $11 r0 *1 16.5,0 res_rppd
R$11 6 46 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $12 r0 *1 18.15,0 res_rppd
R$12 7 46 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $13 r0 *1 19.8,0 res_rppd
R$13 7 47 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $14 r0 *1 21.45,0 res_rppd
R$14 8 47 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $15 r0 *1 23.1,0 res_rppd
R$15 8 48 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $16 r0 *1 24.75,0 res_rppd
R$16 9 48 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $17 r0 *1 26.4,0 res_rppd
R$17 9 49 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $18 r0 *1 28.05,0 res_rppd
R$18 10 49 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $19 r0 *1 29.7,0 res_rppd
R$19 10 50 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $20 r0 *1 31.35,0 res_rppd
R$20 11 50 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $21 r0 *1 33,0 res_rppd
R$21 11 51 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $22 r0 *1 34.65,0 res_rppd
R$22 12 51 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $23 r0 *1 36.3,0 res_rppd
R$23 12 52 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $24 r0 *1 37.95,0 res_rppd
R$24 13 52 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $25 r0 *1 39.6,0 res_rppd
R$25 13 53 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $26 r0 *1 41.25,0 res_rppd
R$26 14 53 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0 ps=0.0 m=1.0
.ENDS sg13g2_RCClampResistor

* Extracted by KLayout with SG13G2 LVS runset on : 03/05/2024 20:22

* cell sg13g2_IOPadInOut16mA
* pin PAD
* pin CORE
* pin sub!
.SUBCKT sg13g2_IOPadInOut16mA PAD CORE sub!
* device instance $1 r0 *1 18.685,171.175 sg13_lv_nmos
M$1 sub! \$84 \$55 sub! sg13_lv_nmos W=3.9299999999999993 L=0.12999999999999998
* device instance $2 r0 *1 19.195,171.175 sg13_lv_nmos
M$2 \$55 \$85 sub! sub! sg13_lv_nmos W=3.9299999999999993 L=0.12999999999999998
* device instance $3 r0 *1 60.255,159.005 sg13_lv_nmos
M$3 \$64 \$66 sub! sub! sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $4 r0 *1 23.485,171.175 sg13_lv_nmos
M$4 sub! \$86 \$85 sub! sg13_lv_nmos W=3.9299999999999993 L=0.12999999999999998
* device instance $5 r0 *1 18.685,159.005 sg13_lv_nmos
M$5 \$54 \$55 sub! sub! sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $6 r0 *1 22.195,159.005 sg13_lv_nmos
M$6 \$56 \$57 sub! sub! sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $7 r0 *1 21.085,171.175 sg13_lv_nmos
M$7 sub! \$84 \$88 sub! sg13_lv_nmos W=3.9299999999999993 L=0.12999999999999998
* device instance $8 r0 *1 21.595,171.175 sg13_lv_nmos
M$8 \$88 \$86 \$57 sub! sg13_lv_nmos W=3.9299999999999993 L=0.12999999999999998
* device instance $9 r0 *1 61.765,159.055 sg13_hv_nmos
M$9 sub! CORE \$66 sub! sg13_hv_nmos W=2.6499999999999995 L=0.4499999999999999
* device instance $10 r0 *1 18.845,155.32 sg13_hv_nmos
M$10 \$48 \$54 sub! sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $11 r0 *1 19.675,155.32 sg13_hv_nmos
M$11 sub! \$55 \$49 sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $12 r0 *1 34.58,10.95 sg13_hv_nmos
M$12 sub! \$6 PAD sub! sg13_hv_nmos W=35.199999999999996 L=0.5999999999999998
* device instance $20 r0 *1 24.525,155.32 sg13_hv_nmos
M$20 sub! \$51 \$32 sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $21 r0 *1 21.015,155.32 sg13_hv_nmos
M$21 sub! \$49 \$6 sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $22 r0 *1 22.355,155.32 sg13_hv_nmos
M$22 \$50 \$56 sub! sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $23 r0 *1 23.185,155.32 sg13_hv_nmos
M$23 sub! \$57 \$51 sub! sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $24 r0 *1 18.685,176.585 sg13_lv_pmos
M$24 \$36 \$84 \$94 \$36 sg13_lv_pmos W=4.409999999999999 L=0.12999999999999995
* device instance $25 r0 *1 19.195,176.585 sg13_lv_pmos
M$25 \$94 \$85 \$55 \$36 sg13_lv_pmos W=4.409999999999999 L=0.12999999999999995
* device instance $26 r0 *1 22.195,163.995 sg13_lv_pmos
M$26 \$56 \$57 \$36 \$36 sg13_lv_pmos W=4.749999999999999 L=0.12999999999999998
* device instance $27 r0 *1 21.085,176.585 sg13_lv_pmos
M$27 \$36 \$84 \$57 \$36 sg13_lv_pmos W=4.409999999999999 L=0.12999999999999995
* device instance $28 r0 *1 21.595,176.585 sg13_lv_pmos
M$28 \$57 \$86 \$36 \$36 sg13_lv_pmos W=4.409999999999999 L=0.12999999999999995
* device instance $29 r0 *1 18.685,163.995 sg13_lv_pmos
M$29 \$54 \$55 \$36 \$36 sg13_lv_pmos W=4.749999999999999 L=0.12999999999999998
* device instance $30 r0 *1 60.255,163.995 sg13_lv_pmos
M$30 \$64 \$66 \$36 \$36 sg13_lv_pmos W=4.749999999999999 L=0.12999999999999998
* device instance $31 r0 *1 23.485,176.585 sg13_lv_pmos
M$31 \$36 \$86 \$85 \$36 sg13_lv_pmos W=4.409999999999999 L=0.12999999999999995
* device instance $32 r0 *1 61.765,163.945 sg13_hv_pmos
M$32 \$36 CORE \$66 \$36 sg13_hv_pmos W=4.6499999999999995 L=0.44999999999999984
* device instance $33 r0 *1 24.525,151.18 sg13_hv_pmos
M$33 \$21 \$51 \$32 \$21 sg13_hv_pmos W=3.899999999999999 L=0.4499999999999999
* device instance $34 r0 *1 21.015,151.18 sg13_hv_pmos
M$34 \$21 \$49 \$6 \$21 sg13_hv_pmos W=3.899999999999999 L=0.4499999999999999
* device instance $35 r0 *1 22.355,151.18 sg13_hv_pmos
M$35 \$50 \$51 \$21 \$21 sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $36 r0 *1 23.185,151.18 sg13_hv_pmos
M$36 \$21 \$50 \$51 \$21 sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $37 r0 *1 18.845,151.18 sg13_hv_pmos
M$37 \$48 \$49 \$21 \$21 sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $38 r0 *1 19.675,151.18 sg13_hv_pmos
M$38 \$21 \$48 \$49 \$21 sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $39 r0 *1 34.58,78.18 sg13_hv_pmos
M$39 \$21 \$32 PAD \$21 sg13_hv_pmos W=106.55999999999996 L=0.5999999999999999
* device instance $55 r0 *1 17.975,12.83 dantenna
D$55 sub! \$6 dantenna A=0.192 P=1.88 m=1
* device instance $56 r0 *1 40,20.44 dantenna
D$56 sub! PAD dantenna A=35.0028 P=58.08 m=2
* device instance $58 r0 *1 65.225,142.54 dantenna
D$58 sub! CORE dantenna A=1.984 P=7.48 m=1
* device instance $59 r0 *1 40,55.96 dpantenna
D$59 PAD \$21 dpantenna A=35.0028 P=58.08 m=2
* device instance $61 r0 *1 17.975,81.19 dpantenna
D$61 \$32 \$21 dpantenna A=0.192 P=1.88 m=1
* device instance $62 r0 *1 63.055,147.51 dpantenna
D$62 CORE \$21 dpantenna A=3.1872 P=11.24 m=1
* device instance $63 r0 *1 60.685,141.11 rppd
R$63 PAD CORE rppd w=1 l=2 ps=0 b=0 m=1
.ENDS sg13g2_IOPadInOut16mA

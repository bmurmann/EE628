* Extracted by KLayout with SG13G2 LVS runset on : 10/05/2024 01:50

* cell Team5
* pin Q
* pin inv_bottom
* pin VDD
* pin nand_B2
* pin Q_N
* pin D
* pin VSS
.SUBCKT Team5 Q inv_bottom VDD nand_B2 Q_N D VSS
* device instance $1 r0 *1 -15.769,-16.292 sg13_lv_nmos
M$1 \$12 \$7 VSS VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $2 r0 *1 -15.259,-16.242 sg13_lv_nmos
M$2 VSS Q \$17 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $3 r0 *1 -14.749,-16.242 sg13_lv_nmos
M$3 \$17 \$42 \$7 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $4 r0 *1 -3.629,-16.242 sg13_lv_nmos
M$4 \$8 \$29 \$15 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $5 r0 *1 -3.119,-16.242 sg13_lv_nmos
M$5 VSS \$14 \$15 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $6 r0 *1 -2.609,-16.292 sg13_lv_nmos
M$6 VSS \$8 \$9 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $7 r0 *1 -36.474,-6.73 sg13_lv_nmos
M$7 \$90 \$42 \$4 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $8 r0 *1 -31.898,-6.73 sg13_lv_nmos
M$8 \$4 \$198 \$47 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $9 r0 *1 -21.672,-10.623 sg13_lv_nmos
M$9 \$19 \$29 \$36 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $10 r0 *1 -20.515,-15.348 sg13_lv_nmos
M$10 \$2 \$12 \$19 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $11 r0 *1 2.137,-15.348 sg13_lv_nmos
M$11 \$2 \$9 \$37 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $12 r0 *1 3.294,-10.623 sg13_lv_nmos
M$12 \$107 \$42 \$37 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $13 r0 *1 13.52,-6.73 sg13_lv_nmos
M$13 \$48 inv_bottom \$5 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $14 r0 *1 18.096,-6.73 sg13_lv_nmos
M$14 \$5 \$29 \$91 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $15 r0 *1 -21.277,-4.14 sg13_lv_nmos
M$15 VSS \$29 \$30 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $16 r0 *1 -17.929,-4.045 sg13_lv_nmos
M$16 VSS Q \$61 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $17 r0 *1 -17.079,-4.14 sg13_lv_nmos
M$17 VSS \$42 \$70 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $18 r0 *1 -16.769,-4.14 sg13_lv_nmos
M$18 \$70 \$61 \$62 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $19 r0 *1 -1.609,-4.14 sg13_lv_nmos
M$19 \$64 \$65 \$69 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $20 r0 *1 -1.299,-4.14 sg13_lv_nmos
M$20 \$69 \$29 VSS VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $21 r0 *1 -0.449,-4.045 sg13_lv_nmos
M$21 VSS \$14 \$65 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $22 r0 *1 2.899,-4.14 sg13_lv_nmos
M$22 \$31 \$42 VSS VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $23 r0 *1 -25.959,1.248 sg13_lv_nmos
M$23 \$47 \$47 VSS VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $24 r0 *1 -25.959,10.794 sg13_lv_nmos
M$24 \$107 \$3 VSS VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $25 r0 *1 7.581,1.248 sg13_lv_nmos
M$25 VSS \$48 \$48 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $26 r0 *1 7.581,10.794 sg13_lv_nmos
M$26 VSS \$6 \$106 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $27 r0 *1 -21.021,13.251 sg13_lv_nmos
M$27 \$107 \$108 \$90 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $28 r0 *1 -16.445,13.251 sg13_lv_nmos
M$28 \$90 \$29 \$3 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $29 r0 *1 -1.933,13.251 sg13_lv_nmos
M$29 \$6 \$42 \$91 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $30 r0 *1 2.643,13.251 sg13_lv_nmos
M$30 \$91 \$108 \$106 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $31 r0 *1 -27.268,20.97 sg13_lv_nmos
M$31 \$134 nand_B2 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $33 r0 *1 -26.238,20.97 sg13_lv_nmos
M$33 \$134 \$199 \$153 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $35 r0 *1 -2.082,20.97 sg13_lv_nmos
M$35 \$141 \$140 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $37 r0 *1 -1.052,20.97 sg13_lv_nmos
M$37 \$141 \$138 \$154 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $39 r0 *1 -24.004,20.995 sg13_lv_nmos
M$39 VSS \$153 \$135 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $43 r0 *1 -20.589,20.995 sg13_lv_nmos
M$43 VSS \$135 \$136 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $47 r0 *1 -17.353,20.995 sg13_lv_nmos
M$47 VSS \$136 \$137 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $51 r0 *1 -13.828,20.995 sg13_lv_nmos
M$51 VSS \$137 \$138 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $55 r0 *1 -9.971,20.995 sg13_lv_nmos
M$55 VSS \$138 inv_bottom VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $59 r0 *1 -6.002,20.995 sg13_lv_nmos
M$59 VSS inv_bottom \$140 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $63 r0 *1 1.602,20.995 sg13_lv_nmos
M$63 VSS \$154 \$142 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $67 r0 *1 4.998,20.995 sg13_lv_nmos
M$67 VSS \$142 \$42 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $75 r0 *1 -33.157,28.963 sg13_lv_nmos
M$75 VSS \$214 nand_B2 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $77 r0 *1 -30.636,28.963 sg13_lv_nmos
M$77 VSS nand_B2 \$216 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $79 r0 *1 -27.99,28.938 sg13_lv_nmos
M$79 \$193 \$216 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $81 r0 *1 -26.96,28.938 sg13_lv_nmos
M$81 \$193 \$140 \$217 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $83 r0 *1 -24.627,28.964 sg13_lv_nmos
M$83 VSS \$217 \$194 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $87 r0 *1 -20.159,28.964 sg13_lv_nmos
M$87 VSS \$194 \$195 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $91 r0 *1 -16.743,28.964 sg13_lv_nmos
M$91 VSS \$195 \$196 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $95 r0 *1 -13.223,28.964 sg13_lv_nmos
M$95 VSS \$196 \$197 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $99 r0 *1 -9.366,28.964 sg13_lv_nmos
M$99 VSS \$197 \$198 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $103 r0 *1 -5.397,28.964 sg13_lv_nmos
M$103 VSS \$198 \$199 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $107 r0 *1 -1.727,28.939 sg13_lv_nmos
M$107 \$200 \$199 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $109 r0 *1 -0.697,28.939 sg13_lv_nmos
M$109 \$200 \$197 \$218 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $111 r0 *1 1.957,28.964 sg13_lv_nmos
M$111 VSS \$218 \$201 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $115 r0 *1 5.353,28.964 sg13_lv_nmos
M$115 VSS \$201 \$29 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $123 r0 *1 -29.808,40.371 sg13_lv_nmos
M$123 VSS \$303 \$326 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $124 r0 *1 -29.808,46.171 sg13_lv_nmos
M$124 VSS \$234 \$347 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $125 r0 *1 -30.676,36.442 sg13_lv_nmos
M$125 VSS \$274 \$14 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $127 r0 *1 -29.656,36.492 sg13_lv_nmos
M$127 VSS D \$274 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $128 r0 *1 -29.766,43.87 sg13_lv_nmos
M$128 D \$360 \$326 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $129 r0 *1 -29.766,49.67 sg13_lv_nmos
M$129 \$360 D \$347 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $130 r0 *1 -27.676,36.262 sg13_lv_nmos
M$130 \$275 D \$285 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $131 r0 *1 -27.366,36.262 sg13_lv_nmos
M$131 \$285 \$262 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $132 r0 *1 -26.786,36.647 sg13_lv_nmos
M$132 VSS \$299 \$263 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $133 r0 *1 -25.696,36.327 sg13_lv_nmos
M$133 VSS \$262 \$287 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $134 r0 *1 -25.386,36.327 sg13_lv_nmos
M$134 \$287 \$263 \$276 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $135 r0 *1 -24.611,37.052 sg13_lv_nmos
M$135 \$275 \$264 \$299 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $136 r0 *1 -24.101,37.052 sg13_lv_nmos
M$136 \$299 \$277 \$276 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $137 r0 *1 -22.841,36.527 sg13_lv_nmos
M$137 VSS \$264 \$277 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $138 r0 *1 -21.741,36.527 sg13_lv_nmos
M$138 VSS \$29 \$264 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $139 r0 *1 -20.531,36.647 sg13_lv_nmos
M$139 \$279 \$264 \$278 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $140 r0 *1 -19.996,36.487 sg13_lv_nmos
M$140 \$263 \$277 \$279 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $141 r0 *1 -18.946,36.262 sg13_lv_nmos
M$141 \$278 \$280 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $142 r0 *1 -18.436,36.262 sg13_lv_nmos
M$142 VSS \$262 \$294 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $143 r0 *1 -18.126,36.262 sg13_lv_nmos
M$143 \$294 \$279 \$280 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $144 r0 *1 -16.086,36.372 sg13_lv_nmos
M$144 VSS \$279 \$266 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $145 r0 *1 -17.106,36.422 sg13_lv_nmos
M$145 VSS \$279 Q_N VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $147 r0 *1 -15.066,36.422 sg13_lv_nmos
M$147 VSS \$266 Q VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $149 r0 *1 -12.295,36.442 sg13_lv_nmos
M$149 VSS \$108 \$262 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $150 r0 *1 -10.86,36.442 sg13_lv_nmos
M$150 VSS \$29 \$281 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $151 r0 *1 -10.307,41.053 sg13_lv_nmos
M$151 \$267 \$29 \$106 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $152 r0 *1 0.059,35.671 sg13_lv_nmos
M$152 VSS \$267 \$233 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $153 r0 *1 0.059,41.332 sg13_lv_nmos
M$153 VSS \$48 \$304 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $154 r0 *1 3.419,42.999 sg13_lv_nmos
M$154 \$303 \$234 \$333 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $155 r0 *1 3.419,37.338 sg13_lv_nmos
M$155 \$234 \$303 \$282 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $156 r0 *1 5.064,37.338 sg13_lv_nmos
M$156 \$282 \$42 \$233 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $157 r0 *1 5.064,42.999 sg13_lv_nmos
M$157 \$333 \$42 \$304 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $158 r0 *1 -15.769,-14.742 sg13_lv_pmos
M$158 \$12 \$7 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $159 r0 *1 -15.259,-14.602 sg13_lv_pmos
M$159 VDD Q \$7 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $160 r0 *1 -14.749,-14.602 sg13_lv_pmos
M$160 \$7 \$42 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $161 r0 *1 -3.629,-14.602 sg13_lv_pmos
M$161 VDD \$29 \$8 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $162 r0 *1 -3.119,-14.602 sg13_lv_pmos
M$162 VDD \$14 \$8 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $163 r0 *1 -2.609,-14.742 sg13_lv_pmos
M$163 VDD \$8 \$9 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $164 r0 *1 -16.04,-10.621 sg13_lv_pmos
M$164 \$19 \$30 \$36 \$26 sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $168 r0 *1 -3.868,-10.621 sg13_lv_pmos
M$168 \$37 \$31 \$107 \$26 sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $172 r0 *1 -17.929,-2.62 sg13_lv_pmos
M$172 \$61 Q VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $173 r0 *1 -17.389,-2.48 sg13_lv_pmos
M$173 VDD \$42 \$62 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $174 r0 *1 -16.879,-2.48 sg13_lv_pmos
M$174 \$62 \$61 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $175 r0 *1 -13.818,-2.992 sg13_lv_pmos
M$175 \$63 \$62 \$19 \$26 sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $176 r0 *1 -4.56,-2.992 sg13_lv_pmos
M$176 \$37 \$64 \$63 \$26 sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $177 r0 *1 -0.449,-2.62 sg13_lv_pmos
M$177 VDD \$14 \$65 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $178 r0 *1 -1.499,-2.48 sg13_lv_pmos
M$178 VDD \$65 \$64 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $179 r0 *1 -0.989,-2.48 sg13_lv_pmos
M$179 \$64 \$29 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $180 r0 *1 -38.017,1.264 sg13_lv_pmos
M$180 \$47 \$47 \$26 \$26 sg13_lv_pmos W=10.0 L=1.5
* device instance $184 r0 *1 -21.267,-2.465 sg13_lv_pmos
M$184 VDD \$29 \$30 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $185 r0 *1 2.889,-2.465 sg13_lv_pmos
M$185 \$31 \$42 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $186 r0 *1 13.999,1.264 sg13_lv_pmos
M$186 \$48 \$48 \$26 \$26 sg13_lv_pmos W=10.0 L=1.5
* device instance $190 r0 *1 -38.017,10.81 sg13_lv_pmos
M$190 \$107 \$3 \$26 \$26 sg13_lv_pmos W=10.0 L=1.5
* device instance $194 r0 *1 13.999,10.81 sg13_lv_pmos
M$194 \$106 \$6 \$26 \$26 sg13_lv_pmos W=10.0 L=1.5
* device instance $198 r0 *1 -27.268,22.655 sg13_lv_pmos
M$198 VDD nand_B2 \$153 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $200 r0 *1 -26.238,22.655 sg13_lv_pmos
M$200 VDD \$199 \$153 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $202 r0 *1 -24.004,22.655 sg13_lv_pmos
M$202 VDD \$153 \$135 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $206 r0 *1 -20.589,22.655 sg13_lv_pmos
M$206 VDD \$135 \$136 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $210 r0 *1 -17.353,22.655 sg13_lv_pmos
M$210 VDD \$136 \$137 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $214 r0 *1 -13.828,22.655 sg13_lv_pmos
M$214 VDD \$137 \$138 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $218 r0 *1 -9.971,22.655 sg13_lv_pmos
M$218 VDD \$138 inv_bottom VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $222 r0 *1 -6.002,22.655 sg13_lv_pmos
M$222 VDD inv_bottom \$140 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $226 r0 *1 -2.082,22.655 sg13_lv_pmos
M$226 VDD \$140 \$154 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $228 r0 *1 -1.052,22.655 sg13_lv_pmos
M$228 VDD \$138 \$154 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $230 r0 *1 1.602,22.655 sg13_lv_pmos
M$230 VDD \$154 \$142 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $234 r0 *1 4.998,22.655 sg13_lv_pmos
M$234 VDD \$142 \$42 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $242 r0 *1 -33.167,30.623 sg13_lv_pmos
M$242 VDD \$214 nand_B2 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $244 r0 *1 -30.646,30.623 sg13_lv_pmos
M$244 VDD nand_B2 \$216 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $246 r0 *1 -27.99,30.623 sg13_lv_pmos
M$246 VDD \$216 \$217 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $248 r0 *1 -26.96,30.623 sg13_lv_pmos
M$248 VDD \$140 \$217 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $250 r0 *1 -24.627,30.624 sg13_lv_pmos
M$250 VDD \$217 \$194 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $254 r0 *1 -20.159,30.624 sg13_lv_pmos
M$254 VDD \$194 \$195 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $258 r0 *1 -16.743,30.624 sg13_lv_pmos
M$258 VDD \$195 \$196 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $262 r0 *1 -13.223,30.624 sg13_lv_pmos
M$262 VDD \$196 \$197 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $266 r0 *1 -9.366,30.624 sg13_lv_pmos
M$266 VDD \$197 \$198 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $270 r0 *1 -5.397,30.624 sg13_lv_pmos
M$270 VDD \$198 \$199 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $274 r0 *1 -1.727,30.624 sg13_lv_pmos
M$274 VDD \$199 \$218 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $276 r0 *1 -0.697,30.624 sg13_lv_pmos
M$276 VDD \$197 \$218 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $278 r0 *1 1.957,30.624 sg13_lv_pmos
M$278 VDD \$218 \$201 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $282 r0 *1 5.353,30.624 sg13_lv_pmos
M$282 VDD \$201 \$29 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $290 r0 *1 -31.066,49.035 sg13_lv_pmos
M$290 \$360 \$234 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $291 r0 *1 -31.066,43.235 sg13_lv_pmos
M$291 D \$303 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $292 r0 *1 -29.656,38.117 sg13_lv_pmos
M$292 VDD D \$274 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $293 r0 *1 -30.676,38.102 sg13_lv_pmos
M$293 VDD \$274 \$14 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $295 r0 *1 -27.786,37.852 sg13_lv_pmos
M$295 VDD D \$275 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $296 r0 *1 -27.276,37.852 sg13_lv_pmos
M$296 VDD \$262 \$275 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $297 r0 *1 -26.826,38.142 sg13_lv_pmos
M$297 VDD \$299 \$263 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $298 r0 *1 -27.624,43.235 sg13_lv_pmos
M$298 VDD \$360 D VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $299 r0 *1 -27.624,49.035 sg13_lv_pmos
M$299 VDD D \$360 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $300 r0 *1 -25.776,38.217 sg13_lv_pmos
M$300 \$299 \$262 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $301 r0 *1 -25.041,38.217 sg13_lv_pmos
M$301 VDD \$263 \$309 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $302 r0 *1 -24.651,38.217 sg13_lv_pmos
M$302 \$309 \$264 \$299 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $303 r0 *1 -24.141,38.217 sg13_lv_pmos
M$303 \$299 \$277 \$275 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $304 r0 *1 -22.441,38.092 sg13_lv_pmos
M$304 \$277 \$264 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $305 r0 *1 -21.716,38.092 sg13_lv_pmos
M$305 VDD \$29 \$264 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $306 r0 *1 -19.586,37.837 sg13_lv_pmos
M$306 \$279 \$277 \$313 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $307 r0 *1 -19.206,37.837 sg13_lv_pmos
M$307 \$313 \$280 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $308 r0 *1 -18.596,37.837 sg13_lv_pmos
M$308 VDD \$262 \$280 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $309 r0 *1 -18.086,37.837 sg13_lv_pmos
M$309 VDD \$279 \$280 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $310 r0 *1 -16.526,37.942 sg13_lv_pmos
M$310 VDD \$279 \$266 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $311 r0 *1 -17.546,38.002 sg13_lv_pmos
M$311 VDD \$279 Q_N VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $313 r0 *1 -20.281,38.127 sg13_lv_pmos
M$313 \$263 \$264 \$279 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $314 r0 *1 -15.441,38.102 sg13_lv_pmos
M$314 VDD \$266 Q VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $316 r0 *1 -12.285,38.117 sg13_lv_pmos
M$316 VDD \$108 \$262 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $317 r0 *1 -10.85,38.117 sg13_lv_pmos
M$317 VDD \$29 \$281 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $318 r0 *1 -9.022,39.053 sg13_lv_pmos
M$318 \$106 \$281 \$267 \$26 sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $319 r0 *1 1.568,42.025 sg13_lv_pmos
M$319 \$26 \$234 \$303 \$26 sg13_lv_pmos W=4.0 L=0.13
* device instance $320 r0 *1 1.568,36.364 sg13_lv_pmos
M$320 \$26 \$303 \$234 \$26 sg13_lv_pmos W=4.0 L=0.13
* device instance $321 r0 *1 6.915,42.025 sg13_lv_pmos
M$321 \$303 \$42 \$26 \$26 sg13_lv_pmos W=4.0 L=0.13
* device instance $322 r0 *1 6.915,36.364 sg13_lv_pmos
M$322 \$234 \$42 \$26 \$26 sg13_lv_pmos W=4.0 L=0.13
* device instance $323 r0 *1 -40.106,-18.735 cap_cmim
C$323 \$3 \$4 cap_cmim w=8.16 l=8.16 m=1
* device instance $324 r0 *1 12.368,-18.735 cap_cmim
C$324 \$6 \$5 cap_cmim w=8.16 l=8.16 m=1
* device instance $325 r0 *1 -30.531,-18.73 cap_cmim
C$325 \$4 \$19 cap_cmim w=5.77 l=5.77 m=1
* device instance $326 r0 *1 -22.287,0.953 cap_cmim
C$326 \$90 \$107 cap_cmim w=8.16 l=8.16 m=1
* device instance $327 r0 *1 5.183,-18.73 cap_cmim
C$327 \$5 \$37 cap_cmim w=5.77 l=5.77 m=1
* device instance $328 r0 *1 -5.451,0.953 cap_cmim
C$328 \$91 \$106 cap_cmim w=8.16 l=8.16 m=1
* device instance $329 r0 *1 -8.533,35.302 cap_cmim
C$329 \$267 VSS cap_cmim w=5.77 l=5.77 m=1
.ENDS Team5

* Extracted by KLayout with SG13G2 LVS runset on : 03/05/2024 20:10

* cell sg13g2_IOPadIOVdd
* pin sub!
.SUBCKT sg13g2_IOPadIOVdd sub!
* device instance $1 r0 *1 8.155,10.95 sg13_hv_nmos
M$1 sub! \$7 \$1 sub! sg13_hv_nmos W=756.7999999999977 L=0.5999999999999998
* device instance $173 r0 *1 3.22,71.54 sg13_hv_nmos
M$173 sub! \$12 \$7 sub! sg13_hv_nmos W=107.99999999999999 L=0.4999999999999999
* device instance $179 r0 *1 13,71.54 sg13_hv_nmos
M$179 sub! \$12 sub! sub! sg13_hv_nmos W=125.99999999999999 L=9.499999999999996
* device instance $199 r0 *1 18.44,94.91 sg13_hv_pmos
M$199 \$1 \$12 \$7 \$1 sg13_hv_pmos W=349.99999999999994 L=0.4999999999999999
* device instance $249 r0 *1 4.765,27.35 dantenna
D$249 sub! \$7 dantenna A=0.192 P=1.88 m=1
* device instance $250 r0 *1 18.875,37.71 rppd
R$250 \$1 \$12 rppd w=1 l=0 ps=0 b=25 m=1
.ENDS sg13g2_IOPadIOVdd

* Extracted by KLayout with SG13G2 LVS runset on : 08/05/2024 07:34

* cell integ_5_splitTop2
* pin sub!
.SUBCKT integ_5_splitTop2 sub!
* device instance $1 r0 *1 -4.307,-17.041 sg13_lv_nmos
M$1 \$7 \$6 \$1 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $2 r0 *1 0.269,-17.041 sg13_lv_nmos
M$2 \$1 \$5 \$8 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $3 r0 *1 -10.246,-9.063 sg13_lv_nmos
M$3 sub! \$7 \$7 sub! sg13_lv_nmos W=2.5 L=1.5
* device instance $4 r0 *1 -10.246,0.483 sg13_lv_nmos
M$4 sub! \$3 \$23 sub! sg13_lv_nmos W=2.5 L=1.5
* device instance $5 r0 *1 -3.828,-9.047 sg13_lv_pmos
M$5 \$7 \$7 \$14 \$14 sg13_lv_pmos W=10.0 L=1.5
* device instance $9 r0 *1 -3.828,0.499 sg13_lv_pmos
M$9 \$23 \$3 \$14 \$14 sg13_lv_pmos W=10.0 L=1.5
* device instance $13 r0 *1 -12.644,-29.041 cap_cmim
C$13 \$1 \$2 cap_cmim w=5.77 l=5.77 m=1
* device instance $14 r0 *1 -5.459,-29.046 cap_cmim
C$14 \$3 \$1 cap_cmim w=8.16 l=8.16 m=1
.ENDS integ_5_splitTop2

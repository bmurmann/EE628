* Extracted by KLayout with SG13G2 LVS runset on : 09/05/2024 23:57

* cell Team5_split2
* pin inv_bottom
* pin VDD
* pin nand_B2
* pin Q_N
* pin Q
* pin D
* pin VSS
.SUBCKT Team5_split2 inv_bottom VDD nand_B2 Q_N Q D VSS
* device instance $1 r0 *1 7.221,-41.489 sg13_lv_nmos
M$1 \$3 nand_B2 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $3 r0 *1 8.251,-41.489 sg13_lv_nmos
M$3 \$3 \$69 \$15 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $5 r0 *1 32.407,-41.489 sg13_lv_nmos
M$5 \$4 \$21 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $7 r0 *1 33.437,-41.489 sg13_lv_nmos
M$7 \$4 \$19 \$22 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $9 r0 *1 10.485,-41.464 sg13_lv_nmos
M$9 VSS \$15 \$16 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $13 r0 *1 13.9,-41.464 sg13_lv_nmos
M$13 VSS \$16 \$17 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $17 r0 *1 17.136,-41.464 sg13_lv_nmos
M$17 VSS \$17 \$18 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $21 r0 *1 20.661,-41.464 sg13_lv_nmos
M$21 VSS \$18 \$19 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $25 r0 *1 24.518,-41.464 sg13_lv_nmos
M$25 VSS \$19 inv_bottom VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $29 r0 *1 28.487,-41.464 sg13_lv_nmos
M$29 VSS inv_bottom \$21 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $33 r0 *1 36.091,-41.464 sg13_lv_nmos
M$33 VSS \$22 \$23 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $37 r0 *1 39.487,-41.464 sg13_lv_nmos
M$37 VSS \$23 \$24 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $45 r0 *1 1.332,-33.496 sg13_lv_nmos
M$45 VSS \$84 nand_B2 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $47 r0 *1 3.853,-33.496 sg13_lv_nmos
M$47 VSS nand_B2 \$86 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $49 r0 *1 6.499,-33.521 sg13_lv_nmos
M$49 \$63 \$86 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $51 r0 *1 7.529,-33.521 sg13_lv_nmos
M$51 \$63 \$21 \$87 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $53 r0 *1 9.862,-33.495 sg13_lv_nmos
M$53 VSS \$87 \$64 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $57 r0 *1 14.33,-33.495 sg13_lv_nmos
M$57 VSS \$64 \$65 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $61 r0 *1 17.746,-33.495 sg13_lv_nmos
M$61 VSS \$65 \$66 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $65 r0 *1 21.266,-33.495 sg13_lv_nmos
M$65 VSS \$66 \$67 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $69 r0 *1 25.123,-33.495 sg13_lv_nmos
M$69 VSS \$67 \$68 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $73 r0 *1 29.092,-33.495 sg13_lv_nmos
M$73 VSS \$68 \$69 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $77 r0 *1 32.762,-33.52 sg13_lv_nmos
M$77 \$70 \$69 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $79 r0 *1 33.792,-33.52 sg13_lv_nmos
M$79 \$70 \$67 \$88 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $81 r0 *1 36.446,-33.495 sg13_lv_nmos
M$81 VSS \$88 \$71 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $85 r0 *1 39.842,-33.495 sg13_lv_nmos
M$85 VSS \$71 \$89 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $93 r0 *1 4.681,-16.288 sg13_lv_nmos
M$93 VSS \$118 \$224 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $94 r0 *1 4.681,-22.088 sg13_lv_nmos
M$94 VSS \$177 \$202 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $95 r0 *1 3.813,-26.017 sg13_lv_nmos
M$95 VSS \$170 \$143 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $97 r0 *1 4.833,-25.967 sg13_lv_nmos
M$97 VSS D \$170 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $98 r0 *1 4.723,-18.589 sg13_lv_nmos
M$98 D \$237 \$202 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $99 r0 *1 4.723,-12.789 sg13_lv_nmos
M$99 \$237 D \$224 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $100 r0 *1 6.813,-26.197 sg13_lv_nmos
M$100 \$144 D \$158 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $101 r0 *1 7.123,-26.197 sg13_lv_nmos
M$101 \$158 \$134 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $102 r0 *1 7.703,-25.812 sg13_lv_nmos
M$102 VSS \$171 \$135 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $103 r0 *1 8.793,-26.132 sg13_lv_nmos
M$103 VSS \$134 \$159 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $104 r0 *1 9.103,-26.132 sg13_lv_nmos
M$104 \$159 \$135 \$145 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $105 r0 *1 9.878,-25.407 sg13_lv_nmos
M$105 \$144 \$136 \$171 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $106 r0 *1 10.388,-25.407 sg13_lv_nmos
M$106 \$171 \$176 \$145 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $107 r0 *1 11.648,-25.932 sg13_lv_nmos
M$107 VSS \$136 \$176 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $108 r0 *1 12.748,-25.932 sg13_lv_nmos
M$108 VSS \$89 \$136 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $109 r0 *1 13.958,-25.812 sg13_lv_nmos
M$109 \$147 \$136 \$146 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $110 r0 *1 14.493,-25.972 sg13_lv_nmos
M$110 \$135 \$176 \$147 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $111 r0 *1 15.543,-26.197 sg13_lv_nmos
M$111 \$146 \$148 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $112 r0 *1 16.053,-26.197 sg13_lv_nmos
M$112 VSS \$134 \$167 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $113 r0 *1 16.363,-26.197 sg13_lv_nmos
M$113 \$167 \$147 \$148 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $114 r0 *1 18.403,-26.087 sg13_lv_nmos
M$114 VSS \$147 \$150 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $115 r0 *1 17.383,-26.037 sg13_lv_nmos
M$115 VSS \$147 Q_N VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $117 r0 *1 19.423,-26.037 sg13_lv_nmos
M$117 VSS \$150 Q VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $119 r0 *1 22.194,-26.017 sg13_lv_nmos
M$119 VSS \$172 \$134 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $120 r0 *1 23.629,-26.017 sg13_lv_nmos
M$120 VSS \$89 \$152 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $121 r0 *1 24.182,-21.406 sg13_lv_nmos
M$121 \$154 \$89 \$153 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $122 r0 *1 34.548,-21.127 sg13_lv_nmos
M$122 VSS \$213 \$188 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $123 r0 *1 34.548,-26.788 sg13_lv_nmos
M$123 VSS \$154 \$117 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $124 r0 *1 37.908,-25.121 sg13_lv_nmos
M$124 \$118 \$177 \$155 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $125 r0 *1 37.908,-19.46 sg13_lv_nmos
M$125 \$177 \$118 \$214 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $126 r0 *1 39.553,-25.121 sg13_lv_nmos
M$126 \$155 \$24 \$117 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $127 r0 *1 39.553,-19.46 sg13_lv_nmos
M$127 \$214 \$24 \$188 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $128 r0 *1 7.221,-39.804 sg13_lv_pmos
M$128 VDD nand_B2 \$15 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $130 r0 *1 8.251,-39.804 sg13_lv_pmos
M$130 VDD \$69 \$15 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $132 r0 *1 10.485,-39.804 sg13_lv_pmos
M$132 VDD \$15 \$16 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $136 r0 *1 13.9,-39.804 sg13_lv_pmos
M$136 VDD \$16 \$17 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $140 r0 *1 17.136,-39.804 sg13_lv_pmos
M$140 VDD \$17 \$18 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $144 r0 *1 20.661,-39.804 sg13_lv_pmos
M$144 VDD \$18 \$19 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $148 r0 *1 24.518,-39.804 sg13_lv_pmos
M$148 VDD \$19 inv_bottom VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $152 r0 *1 28.487,-39.804 sg13_lv_pmos
M$152 VDD inv_bottom \$21 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $156 r0 *1 32.407,-39.804 sg13_lv_pmos
M$156 VDD \$21 \$22 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $158 r0 *1 33.437,-39.804 sg13_lv_pmos
M$158 VDD \$19 \$22 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $160 r0 *1 36.091,-39.804 sg13_lv_pmos
M$160 VDD \$22 \$23 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $164 r0 *1 39.487,-39.804 sg13_lv_pmos
M$164 VDD \$23 \$24 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $172 r0 *1 1.322,-31.836 sg13_lv_pmos
M$172 VDD \$84 nand_B2 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $174 r0 *1 3.843,-31.836 sg13_lv_pmos
M$174 VDD nand_B2 \$86 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $176 r0 *1 6.499,-31.836 sg13_lv_pmos
M$176 VDD \$86 \$87 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $178 r0 *1 7.529,-31.836 sg13_lv_pmos
M$178 VDD \$21 \$87 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $180 r0 *1 9.862,-31.835 sg13_lv_pmos
M$180 VDD \$87 \$64 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $184 r0 *1 14.33,-31.835 sg13_lv_pmos
M$184 VDD \$64 \$65 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $188 r0 *1 17.746,-31.835 sg13_lv_pmos
M$188 VDD \$65 \$66 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $192 r0 *1 21.266,-31.835 sg13_lv_pmos
M$192 VDD \$66 \$67 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $196 r0 *1 25.123,-31.835 sg13_lv_pmos
M$196 VDD \$67 \$68 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $200 r0 *1 29.092,-31.835 sg13_lv_pmos
M$200 VDD \$68 \$69 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $204 r0 *1 32.762,-31.835 sg13_lv_pmos
M$204 VDD \$69 \$88 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $206 r0 *1 33.792,-31.835 sg13_lv_pmos
M$206 VDD \$67 \$88 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $208 r0 *1 36.446,-31.835 sg13_lv_pmos
M$208 VDD \$88 \$71 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $212 r0 *1 39.842,-31.835 sg13_lv_pmos
M$212 VDD \$71 \$89 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $220 r0 *1 3.423,-13.424 sg13_lv_pmos
M$220 \$237 \$118 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $221 r0 *1 3.423,-19.224 sg13_lv_pmos
M$221 D \$177 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $222 r0 *1 4.833,-24.342 sg13_lv_pmos
M$222 VDD D \$170 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $223 r0 *1 3.813,-24.357 sg13_lv_pmos
M$223 VDD \$170 \$143 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $225 r0 *1 6.703,-24.607 sg13_lv_pmos
M$225 VDD D \$144 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $226 r0 *1 7.213,-24.607 sg13_lv_pmos
M$226 VDD \$134 \$144 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $227 r0 *1 7.663,-24.317 sg13_lv_pmos
M$227 VDD \$171 \$135 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $228 r0 *1 6.865,-13.424 sg13_lv_pmos
M$228 VDD D \$237 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $229 r0 *1 6.865,-19.224 sg13_lv_pmos
M$229 VDD \$237 D VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $230 r0 *1 8.713,-24.242 sg13_lv_pmos
M$230 \$171 \$134 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $231 r0 *1 9.448,-24.242 sg13_lv_pmos
M$231 VDD \$135 \$181 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $232 r0 *1 9.838,-24.242 sg13_lv_pmos
M$232 \$181 \$136 \$171 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $233 r0 *1 10.348,-24.242 sg13_lv_pmos
M$233 \$171 \$176 \$144 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $234 r0 *1 12.048,-24.367 sg13_lv_pmos
M$234 \$176 \$136 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $235 r0 *1 12.773,-24.367 sg13_lv_pmos
M$235 VDD \$89 \$136 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $236 r0 *1 14.903,-24.622 sg13_lv_pmos
M$236 \$147 \$176 \$184 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $237 r0 *1 15.283,-24.622 sg13_lv_pmos
M$237 \$184 \$148 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $238 r0 *1 15.893,-24.622 sg13_lv_pmos
M$238 VDD \$134 \$148 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $239 r0 *1 16.403,-24.622 sg13_lv_pmos
M$239 VDD \$147 \$148 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $240 r0 *1 17.963,-24.517 sg13_lv_pmos
M$240 VDD \$147 \$150 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $241 r0 *1 16.943,-24.457 sg13_lv_pmos
M$241 VDD \$147 Q_N VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $243 r0 *1 14.208,-24.332 sg13_lv_pmos
M$243 \$135 \$136 \$147 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $244 r0 *1 19.048,-24.357 sg13_lv_pmos
M$244 VDD \$150 Q VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $246 r0 *1 22.204,-24.342 sg13_lv_pmos
M$246 VDD \$172 \$134 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $247 r0 *1 23.639,-24.342 sg13_lv_pmos
M$247 VDD \$89 \$152 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $248 r0 *1 25.467,-23.406 sg13_lv_pmos
M$248 \$153 \$152 \$154 \$116 sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $249 r0 *1 36.057,-26.095 sg13_lv_pmos
M$249 \$116 \$177 \$118 \$116 sg13_lv_pmos W=4.0 L=0.13
* device instance $250 r0 *1 36.057,-20.434 sg13_lv_pmos
M$250 \$116 \$118 \$177 \$116 sg13_lv_pmos W=4.0 L=0.13
* device instance $251 r0 *1 41.404,-20.434 sg13_lv_pmos
M$251 \$177 \$24 \$116 \$116 sg13_lv_pmos W=4.0 L=0.13
* device instance $252 r0 *1 41.404,-26.095 sg13_lv_pmos
M$252 \$118 \$24 \$116 \$116 sg13_lv_pmos W=4.0 L=0.13
* device instance $253 r0 *1 25.956,-27.157 cap_cmim
C$253 \$154 VSS cap_cmim w=5.77 l=5.77 m=1
.ENDS Team5_split2

* Extracted by KLayout with SG13G2 LVS runset on : 29/04/2024 21:56

* cell sg13g2_Clamp_P20N0D
.SUBCKT sg13g2_Clamp_P20N0D
* device instance $1 r0 *1 25.52,13.18 sg13_hv_pmos
M$1 iovdd \$6 pad iovdd sg13_hv_pmos W=266.3999999999999 L=0.5999999999999999
* device instance $41 r0 *1 66.305,2.75 res_rppd
R$41 iovdd \$6 res_rppd w=0.4999999999999999 l=12.899999999999997 b=0.0 ps=0.0
+ m=1.0
.ENDS sg13g2_Clamp_P20N0D

* Extracted by KLayout with SG13G2 LVS runset on : 05/05/2024 00:53

* cell Team3
* pin sub!
.SUBCKT Team3 sub!
* device instance $1 r0 *1 19.83,1.155 sg13_lv_nmos
M$1 \$4 \$47 sub! sub! sg13_lv_nmos W=1.4399999999999997 L=0.12999999999999998
* device instance $3 r0 *1 20.86,1.155 sg13_lv_nmos
M$3 \$4 \$3 \$5 sub! sg13_lv_nmos W=1.4399999999999997 L=0.12999999999999998
* device instance $5 r0 *1 39.99,1.155 sg13_lv_nmos
M$5 \$12 \$11 sub! sub! sg13_lv_nmos W=1.4399999999999997 L=0.12999999999999998
* device instance $7 r0 *1 41.02,1.155 sg13_lv_nmos
M$7 \$12 \$9 \$13 sub! sg13_lv_nmos W=1.4399999999999997 L=0.12999999999999998
* device instance $9 r0 *1 22.635,1.18 sg13_lv_nmos
M$9 sub! \$5 \$6 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $13 r0 *1 25.515,1.18 sg13_lv_nmos
M$13 sub! \$6 \$7 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $17 r0 *1 28.395,1.18 sg13_lv_nmos
M$17 sub! \$7 \$8 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $21 r0 *1 31.275,1.18 sg13_lv_nmos
M$21 sub! \$8 \$9 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $25 r0 *1 34.155,1.18 sg13_lv_nmos
M$25 sub! \$9 \$10 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $29 r0 *1 37.035,1.18 sg13_lv_nmos
M$29 sub! \$10 \$11 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $33 r0 *1 42.795,1.18 sg13_lv_nmos
M$33 sub! \$13 \$14 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $37 r0 *1 45.615,1.18 sg13_lv_nmos
M$37 sub! \$14 \$15 sub! sg13_lv_nmos W=5.92 L=0.12999999999999995
* device instance $45 r0 *1 15.935,6.98 sg13_lv_nmos
M$45 sub! \$64 \$3 sub! sg13_lv_nmos W=1.4799999999999998 L=0.12999999999999995
* device instance $47 r0 *1 17.855,6.98 sg13_lv_nmos
M$47 sub! \$3 \$39 sub! sg13_lv_nmos W=1.4799999999999998 L=0.12999999999999995
* device instance $49 r0 *1 19.83,6.955 sg13_lv_nmos
M$49 \$40 \$11 sub! sub! sg13_lv_nmos W=1.4399999999999997 L=0.12999999999999998
* device instance $51 r0 *1 20.86,6.955 sg13_lv_nmos
M$51 \$40 \$39 \$41 sub! sg13_lv_nmos W=1.4399999999999997 L=0.12999999999999998
* device instance $53 r0 *1 22.635,6.98 sg13_lv_nmos
M$53 sub! \$41 \$42 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $57 r0 *1 25.515,6.98 sg13_lv_nmos
M$57 sub! \$42 \$43 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $61 r0 *1 28.395,6.98 sg13_lv_nmos
M$61 sub! \$43 \$44 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $65 r0 *1 31.275,6.98 sg13_lv_nmos
M$65 sub! \$44 \$45 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $69 r0 *1 34.155,6.98 sg13_lv_nmos
M$69 sub! \$45 \$46 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $73 r0 *1 37.035,6.98 sg13_lv_nmos
M$73 sub! \$46 \$47 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $77 r0 *1 39.99,6.955 sg13_lv_nmos
M$77 \$48 \$47 sub! sub! sg13_lv_nmos W=1.4399999999999997 L=0.12999999999999998
* device instance $79 r0 *1 41.02,6.955 sg13_lv_nmos
M$79 \$48 \$45 \$49 sub! sg13_lv_nmos W=1.4399999999999997 L=0.12999999999999998
* device instance $81 r0 *1 42.795,6.98 sg13_lv_nmos
M$81 sub! \$49 \$50 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $85 r0 *1 45.615,6.98 sg13_lv_nmos
M$85 sub! \$50 \$51 sub! sg13_lv_nmos W=5.92 L=0.12999999999999995
* device instance $93 r0 *1 3.27,20.415 sg13_lv_nmos
M$93 sub! \$51 \$88 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $94 r0 *1 4.36,20.51 sg13_lv_nmos
M$94 sub! \$65 \$89 sub! sg13_lv_nmos W=0.5499999999999999 L=0.12999999999999995
* device instance $95 r0 *1 5.21,20.415 sg13_lv_nmos
M$95 sub! \$15 \$103 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $96 r0 *1 5.52,20.415 sg13_lv_nmos
M$96 \$103 \$89 \$90 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $97 r0 *1 6.85,20.575 sg13_lv_nmos
M$97 \$95 \$15 \$107 sub! sg13_lv_nmos W=0.6399999999999999
+ L=0.12999999999999995
* device instance $98 r0 *1 7.36,20.575 sg13_lv_nmos
M$98 sub! \$65 \$107 sub! sg13_lv_nmos W=0.6399999999999999
+ L=0.12999999999999995
* device instance $99 r0 *1 7.87,20.525 sg13_lv_nmos
M$99 sub! \$95 \$81 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $100 r0 *1 11.655,22.475 sg13_lv_nmos
M$100 \$121 \$81 \$122 sub! sg13_lv_nmos W=0.4999999999999999
+ L=0.12999999999999998
* device instance $101 r0 *1 24.37,20.04 sg13_lv_nmos
M$101 \$82 \$46 \$97 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $102 r0 *1 24.37,20.55 sg13_lv_nmos
M$102 \$97 \$15 \$179 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $103 r0 *1 24.37,21.83 sg13_lv_nmos
M$103 \$211 \$51 \$179 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $104 r0 *1 24.37,22.34 sg13_lv_nmos
M$104 \$179 \$66 \$123 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $105 r0 *1 39.325,20.415 sg13_lv_nmos
M$105 sub! \$15 \$91 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $106 r0 *1 40.415,20.51 sg13_lv_nmos
M$106 sub! \$67 \$92 sub! sg13_lv_nmos W=0.5499999999999999
+ L=0.12999999999999995
* device instance $107 r0 *1 41.265,20.415 sg13_lv_nmos
M$107 sub! \$51 \$114 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $108 r0 *1 41.575,20.415 sg13_lv_nmos
M$108 \$114 \$92 \$93 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $109 r0 *1 42.905,20.575 sg13_lv_nmos
M$109 \$98 \$51 \$110 sub! sg13_lv_nmos W=0.6399999999999999
+ L=0.12999999999999995
* device instance $110 r0 *1 43.415,20.575 sg13_lv_nmos
M$110 sub! \$67 \$110 sub! sg13_lv_nmos W=0.6399999999999999
+ L=0.12999999999999995
* device instance $111 r0 *1 43.925,20.525 sg13_lv_nmos
M$111 sub! \$98 \$83 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $112 r0 *1 47.71,22.475 sg13_lv_nmos
M$112 \$121 \$83 \$124 sub! sg13_lv_nmos W=0.4999999999999999
+ L=0.12999999999999998
* device instance $113 r0 *1 60.425,21.83 sg13_lv_nmos
M$113 \$212 \$15 \$180 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $114 r0 *1 60.425,22.34 sg13_lv_nmos
M$114 \$180 \$66 \$125 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $115 r0 *1 60.425,20.04 sg13_lv_nmos
M$115 \$84 \$10 \$99 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $116 r0 *1 60.425,20.55 sg13_lv_nmos
M$116 \$99 \$51 \$180 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $117 r0 *1 75.425,20.53 sg13_lv_nmos
M$117 sub! \$51 \$94 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $118 r0 *1 90.915,23.83 sg13_lv_nmos
M$118 \$150 \$149 \$168 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $119 r0 *1 91.225,23.83 sg13_lv_nmos
M$119 \$168 \$140 sub! sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $120 r0 *1 91.805,24.215 sg13_lv_nmos
M$120 sub! \$171 \$141 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $121 r0 *1 92.895,23.895 sg13_lv_nmos
M$121 sub! \$140 \$166 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $122 r0 *1 93.205,23.895 sg13_lv_nmos
M$122 \$166 \$141 \$151 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $123 r0 *1 95.75,24.095 sg13_lv_nmos
M$123 sub! \$142 \$181 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $124 r0 *1 96.85,24.095 sg13_lv_nmos
M$124 sub! \$51 \$142 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $125 r0 *1 98.06,24.215 sg13_lv_nmos
M$125 \$153 \$142 \$152 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $126 r0 *1 98.595,24.055 sg13_lv_nmos
M$126 \$141 \$181 \$153 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $127 r0 *1 99.645,23.83 sg13_lv_nmos
M$127 \$152 \$154 sub! sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $128 r0 *1 100.155,23.83 sg13_lv_nmos
M$128 sub! \$140 \$159 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $129 r0 *1 100.465,23.83 sg13_lv_nmos
M$129 \$159 \$153 \$154 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $130 r0 *1 102.505,23.94 sg13_lv_nmos
M$130 sub! \$153 \$144 sub! sg13_lv_nmos W=0.6399999999999999
+ L=0.12999999999999995
* device instance $131 r0 *1 101.485,23.99 sg13_lv_nmos
M$131 sub! \$153 \$143 sub! sg13_lv_nmos W=1.4799999999999998
+ L=0.12999999999999995
* device instance $133 r0 *1 103.525,23.99 sg13_lv_nmos
M$133 sub! \$144 \$65 sub! sg13_lv_nmos W=1.4799999999999998
+ L=0.12999999999999995
* device instance $135 r0 *1 105.21,24.01 sg13_lv_nmos
M$135 sub! \$65 \$126 sub! sg13_lv_nmos W=1.4799999999999998
+ L=0.12999999999999995
* device instance $137 r0 *1 107,24.005 sg13_lv_nmos
M$137 \$140 \$66 sub! sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $138 r0 *1 3.495,25.675 sg13_lv_nmos
M$138 \$169 \$51 \$122 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $139 r0 *1 26.64,27.065 sg13_lv_nmos
M$139 sub! \$211 \$123 sub! sg13_lv_nmos W=2.4999999999999996
+ L=1.4999999999999996
* device instance $140 r0 *1 32.64,27.065 sg13_lv_nmos
M$140 sub! \$82 \$82 sub! sg13_lv_nmos W=2.4999999999999996 L=1.4999999999999996
* device instance $141 r0 *1 39.55,25.675 sg13_lv_nmos
M$141 \$123 \$15 \$124 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $142 r0 *1 62.695,27.065 sg13_lv_nmos
M$142 sub! \$212 \$125 sub! sg13_lv_nmos W=2.4999999999999996
+ L=1.4999999999999996
* device instance $143 r0 *1 68.695,27.065 sg13_lv_nmos
M$143 sub! \$84 \$84 sub! sg13_lv_nmos W=2.4999999999999996 L=1.4999999999999996
* device instance $144 r0 *1 75.05,27.5 sg13_lv_nmos
M$144 \$170 \$51 \$125 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $145 r0 *1 79.96,30.51 sg13_lv_nmos
M$145 sub! \$84 \$216 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.9999999999999998
* device instance $146 r0 *1 84.885,30.51 sg13_lv_nmos
M$146 sub! \$170 \$217 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.9999999999999998
* device instance $147 r0 *1 93.98,24.62 sg13_lv_nmos
M$147 \$150 \$142 \$171 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $148 r0 *1 94.49,24.62 sg13_lv_nmos
M$148 \$171 \$181 \$151 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $149 r0 *1 102.795,29.47 sg13_lv_nmos
M$149 sub! \$213 \$67 sub! sg13_lv_nmos W=1.4799999999999998
+ L=0.12999999999999995
* device instance $151 r0 *1 102.845,30.49 sg13_lv_nmos
M$151 sub! \$149 \$213 sub! sg13_lv_nmos W=0.6399999999999999
+ L=0.12999999999999995
* device instance $152 r0 *1 92.75,31.29 sg13_lv_nmos
M$152 sub! \$235 \$218 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $153 r0 *1 99.69,31.28 sg13_lv_nmos
M$153 sub! \$234 \$219 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $154 r0 *1 79.855,31.99 sg13_lv_nmos
M$154 \$216 \$15 \$228 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $155 r0 *1 84.795,31.99 sg13_lv_nmos
M$155 \$217 \$15 \$229 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $156 r0 *1 93.03,32.795 sg13_lv_nmos
M$156 \$218 \$149 \$236 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $157 r0 *1 99.34,32.76 sg13_lv_nmos
M$157 \$219 \$236 \$149 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $158 r0 *1 79.835,33.77 sg13_lv_nmos
M$158 \$228 \$235 \$234 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $159 r0 *1 84.62,33.77 sg13_lv_nmos
M$159 \$229 \$234 \$235 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $160 r0 *1 19.83,2.84 sg13_lv_pmos
M$160 \$26 \$47 \$5 \$26 sg13_lv_pmos W=2.2399999999999998 L=0.12999999999999995
* device instance $162 r0 *1 20.86,2.84 sg13_lv_pmos
M$162 \$26 \$3 \$5 \$26 sg13_lv_pmos W=2.2399999999999998 L=0.12999999999999995
* device instance $164 r0 *1 22.635,2.84 sg13_lv_pmos
M$164 \$26 \$5 \$6 \$26 sg13_lv_pmos W=4.4799999999999995 L=0.12999999999999995
* device instance $168 r0 *1 25.515,2.84 sg13_lv_pmos
M$168 \$26 \$6 \$7 \$26 sg13_lv_pmos W=4.4799999999999995 L=0.12999999999999995
* device instance $172 r0 *1 28.395,2.84 sg13_lv_pmos
M$172 \$26 \$7 \$8 \$26 sg13_lv_pmos W=4.4799999999999995 L=0.12999999999999995
* device instance $176 r0 *1 31.275,2.84 sg13_lv_pmos
M$176 \$26 \$8 \$9 \$26 sg13_lv_pmos W=4.4799999999999995 L=0.12999999999999995
* device instance $180 r0 *1 34.155,2.84 sg13_lv_pmos
M$180 \$26 \$9 \$10 \$26 sg13_lv_pmos W=4.4799999999999995 L=0.12999999999999995
* device instance $184 r0 *1 37.035,2.84 sg13_lv_pmos
M$184 \$26 \$10 \$11 \$26 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $188 r0 *1 39.99,2.84 sg13_lv_pmos
M$188 \$26 \$11 \$13 \$26 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $190 r0 *1 41.02,2.84 sg13_lv_pmos
M$190 \$26 \$9 \$13 \$26 sg13_lv_pmos W=2.2399999999999998 L=0.12999999999999995
* device instance $192 r0 *1 42.795,2.84 sg13_lv_pmos
M$192 \$26 \$13 \$14 \$26 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $196 r0 *1 45.615,2.84 sg13_lv_pmos
M$196 \$26 \$14 \$15 \$26 sg13_lv_pmos W=8.959999999999999 L=0.12999999999999995
* device instance $204 r0 *1 15.925,8.64 sg13_lv_pmos
M$204 \$26 \$64 \$3 \$26 sg13_lv_pmos W=2.2399999999999998 L=0.12999999999999995
* device instance $206 r0 *1 17.845,8.64 sg13_lv_pmos
M$206 \$26 \$3 \$39 \$26 sg13_lv_pmos W=2.2399999999999998 L=0.12999999999999995
* device instance $208 r0 *1 19.83,8.64 sg13_lv_pmos
M$208 \$26 \$11 \$41 \$26 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $210 r0 *1 20.86,8.64 sg13_lv_pmos
M$210 \$26 \$39 \$41 \$26 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $212 r0 *1 22.635,8.64 sg13_lv_pmos
M$212 \$26 \$41 \$42 \$26 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $216 r0 *1 25.515,8.64 sg13_lv_pmos
M$216 \$26 \$42 \$43 \$26 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $220 r0 *1 28.395,8.64 sg13_lv_pmos
M$220 \$26 \$43 \$44 \$26 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $224 r0 *1 31.275,8.64 sg13_lv_pmos
M$224 \$26 \$44 \$45 \$26 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $228 r0 *1 34.155,8.64 sg13_lv_pmos
M$228 \$26 \$45 \$46 \$26 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $232 r0 *1 37.035,8.64 sg13_lv_pmos
M$232 \$26 \$46 \$47 \$26 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $236 r0 *1 39.99,8.64 sg13_lv_pmos
M$236 \$26 \$47 \$49 \$26 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $238 r0 *1 41.02,8.64 sg13_lv_pmos
M$238 \$26 \$45 \$49 \$26 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $240 r0 *1 42.795,8.64 sg13_lv_pmos
M$240 \$26 \$49 \$50 \$26 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $244 r0 *1 45.615,8.64 sg13_lv_pmos
M$244 \$26 \$50 \$51 \$26 sg13_lv_pmos W=8.959999999999999 L=0.12999999999999995
* device instance $252 r0 *1 3.28,22.09 sg13_lv_pmos
M$252 \$26 \$51 \$88 \$26 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $253 r0 *1 4.36,21.935 sg13_lv_pmos
M$253 \$89 \$65 \$26 \$26 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $254 r0 *1 4.9,22.075 sg13_lv_pmos
M$254 \$26 \$15 \$90 \$26 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $255 r0 *1 5.41,22.075 sg13_lv_pmos
M$255 \$90 \$89 \$26 \$26 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $256 r0 *1 4.995,25.675 sg13_lv_pmos
M$256 \$169 \$88 \$122 \$215 sg13_lv_pmos W=5.999999999999998
+ L=0.12999999999999998
* device instance $259 r0 *1 6.85,22.215 sg13_lv_pmos
M$259 \$26 \$15 \$95 \$26 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $260 r0 *1 7.36,22.215 sg13_lv_pmos
M$260 \$26 \$65 \$95 \$26 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $261 r0 *1 7.87,22.075 sg13_lv_pmos
M$261 \$26 \$95 \$81 \$26 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $262 r0 *1 9.97,21.765 sg13_lv_pmos
M$262 \$96 \$90 \$122 \$215 sg13_lv_pmos W=1.4999999999999998
+ L=0.12999999999999995
* device instance $263 r0 *1 39.335,22.09 sg13_lv_pmos
M$263 \$26 \$15 \$91 \$26 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $264 r0 *1 40.415,21.935 sg13_lv_pmos
M$264 \$92 \$67 \$26 \$26 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $265 r0 *1 40.955,22.075 sg13_lv_pmos
M$265 \$26 \$51 \$93 \$26 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $266 r0 *1 41.465,22.075 sg13_lv_pmos
M$266 \$93 \$92 \$26 \$26 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $267 r0 *1 41.05,25.675 sg13_lv_pmos
M$267 \$123 \$91 \$124 \$215 sg13_lv_pmos W=5.999999999999998
+ L=0.12999999999999998
* device instance $270 r0 *1 42.905,22.215 sg13_lv_pmos
M$270 \$26 \$51 \$98 \$26 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $271 r0 *1 43.415,22.215 sg13_lv_pmos
M$271 \$26 \$67 \$98 \$26 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $272 r0 *1 43.925,22.075 sg13_lv_pmos
M$272 \$26 \$98 \$83 \$26 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $273 r0 *1 46.025,21.765 sg13_lv_pmos
M$273 \$96 \$93 \$124 \$215 sg13_lv_pmos W=1.4999999999999998
+ L=0.12999999999999995
* device instance $274 r0 *1 75.15,25.115 sg13_lv_pmos
M$274 \$170 \$94 \$125 \$215 sg13_lv_pmos W=5.999999999999998
+ L=0.12999999999999998
* device instance $277 r0 *1 75.435,22.205 sg13_lv_pmos
M$277 \$26 \$51 \$94 \$26 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $278 r0 *1 90.805,25.42 sg13_lv_pmos
M$278 \$26 \$149 \$150 \$26 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $279 r0 *1 91.315,25.42 sg13_lv_pmos
M$279 \$26 \$140 \$150 \$26 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $280 r0 *1 91.765,25.71 sg13_lv_pmos
M$280 \$26 \$171 \$141 \$26 sg13_lv_pmos W=0.9999999999999998
+ L=0.12999999999999998
* device instance $281 r0 *1 92.815,25.785 sg13_lv_pmos
M$281 \$171 \$140 \$26 \$26 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $282 r0 *1 93.55,25.785 sg13_lv_pmos
M$282 \$26 \$141 \$204 \$26 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $283 r0 *1 93.94,25.785 sg13_lv_pmos
M$283 \$204 \$142 \$171 \$26 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $284 r0 *1 94.45,25.785 sg13_lv_pmos
M$284 \$171 \$181 \$150 \$26 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $285 r0 *1 96.15,25.66 sg13_lv_pmos
M$285 \$181 \$142 \$26 \$26 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $286 r0 *1 96.875,25.66 sg13_lv_pmos
M$286 \$26 \$51 \$142 \$26 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $287 r0 *1 99.005,25.405 sg13_lv_pmos
M$287 \$153 \$181 \$184 \$26 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $288 r0 *1 99.385,25.405 sg13_lv_pmos
M$288 \$184 \$154 \$26 \$26 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $289 r0 *1 99.995,25.405 sg13_lv_pmos
M$289 \$26 \$140 \$154 \$26 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $290 r0 *1 100.505,25.405 sg13_lv_pmos
M$290 \$26 \$153 \$154 \$26 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $291 r0 *1 102.065,25.51 sg13_lv_pmos
M$291 \$26 \$153 \$144 \$26 sg13_lv_pmos W=0.9999999999999998
+ L=0.12999999999999998
* device instance $292 r0 *1 101.045,25.57 sg13_lv_pmos
M$292 \$26 \$153 \$143 \$26 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $294 r0 *1 98.31,25.695 sg13_lv_pmos
M$294 \$141 \$142 \$153 \$26 sg13_lv_pmos W=0.9999999999999998
+ L=0.12999999999999998
* device instance $295 r0 *1 103.15,25.67 sg13_lv_pmos
M$295 \$26 \$144 \$65 \$26 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $297 r0 *1 105.2,25.67 sg13_lv_pmos
M$297 \$26 \$65 \$126 \$26 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $299 r0 *1 106.99,25.68 sg13_lv_pmos
M$299 \$140 \$66 \$26 \$26 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $300 r0 *1 26.64,29.975 sg13_lv_pmos
M$300 \$123 \$211 \$215 \$215 sg13_lv_pmos W=9.999999999999998
+ L=1.4999999999999996
* device instance $304 r0 *1 32.64,29.975 sg13_lv_pmos
M$304 \$82 \$82 \$215 \$215 sg13_lv_pmos W=9.999999999999998
+ L=1.4999999999999996
* device instance $308 r0 *1 62.695,29.975 sg13_lv_pmos
M$308 \$125 \$212 \$215 \$215 sg13_lv_pmos W=9.999999999999998
+ L=1.4999999999999996
* device instance $312 r0 *1 68.695,29.975 sg13_lv_pmos
M$312 \$84 \$84 \$215 \$215 sg13_lv_pmos W=9.999999999999998
+ L=1.4999999999999996
* device instance $316 r0 *1 78.41,37.315 sg13_lv_pmos
M$316 \$215 \$15 \$234 \$215 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $317 r0 *1 81.055,37.315 sg13_lv_pmos
M$317 \$234 \$235 \$215 \$215 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $318 r0 *1 83.41,37.315 sg13_lv_pmos
M$318 \$215 \$234 \$235 \$215 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $319 r0 *1 86.045,37.315 sg13_lv_pmos
M$319 \$235 \$15 \$215 \$215 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $320 r0 *1 91.51,36.615 sg13_lv_pmos
M$320 \$26 \$235 \$236 \$26 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $321 r0 *1 94.18,36.615 sg13_lv_pmos
M$321 \$236 \$149 \$26 \$26 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $322 r0 *1 98.19,36.615 sg13_lv_pmos
M$322 \$26 \$236 \$149 \$26 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $323 r0 *1 100.86,36.615 sg13_lv_pmos
M$323 \$149 \$234 \$26 \$26 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $324 r0 *1 104.455,29.47 sg13_lv_pmos
M$324 \$26 \$213 \$67 \$26 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $326 r0 *1 104.47,30.49 sg13_lv_pmos
M$326 \$26 \$149 \$213 \$26 sg13_lv_pmos W=0.9999999999999998
+ L=0.12999999999999998
* device instance $327 r0 *1 79.38,19.465 cap_cmim
C$327 \$170 sub! cap_cmim w=5.77 l=5.77 m=1
* device instance $328 r0 *1 49.935,19.55 cap_cmim
C$328 \$99 \$124 cap_cmim w=5.77 l=5.77 m=1
* device instance $329 r0 *1 0.19,28.19 cap_cmim
C$329 \$179 \$123 cap_cmim w=8.16 l=8.16 m=1
* device instance $330 r0 *1 13.88,19.55 cap_cmim
C$330 \$97 \$122 cap_cmim w=5.77 l=5.77 m=1
* device instance $331 r0 *1 36.245,28.19 cap_cmim
C$331 \$180 \$125 cap_cmim w=8.16 l=8.16 m=1
* device instance $332 r0 *1 11.11,29.165 cap_cmim
C$332 \$211 \$97 cap_cmim w=8.16 l=8.16 m=1
* device instance $333 r0 *1 47.165,29.165 cap_cmim
C$333 \$212 \$99 cap_cmim w=8.16 l=8.16 m=1
.ENDS Team3

* Extracted by KLayout with SG13G2 LVS runset on : 09/05/2024 08:22

* cell comp_5_split1
* pin sub!
.SUBCKT comp_5_split1 sub!
* device instance $1 r0 *1 1.661,-3.011 sg13_lv_nmos
M$1 \$5 \$2 \$6 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $2 r0 *1 3.306,-3.011 sg13_lv_nmos
M$2 \$6 \$3 \$7 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $3 r0 *1 6.666,-1.344 sg13_lv_nmos
M$3 \$5 \$12 sub! sub! sg13_lv_nmos W=2.0 L=1.0
* device instance $4 r0 *1 -0.19,-2.037 sg13_lv_pmos
M$4 \$4 \$2 \$7 \$4 sg13_lv_pmos W=4.0 L=0.13
* device instance $5 r0 *1 5.157,-2.037 sg13_lv_pmos
M$5 \$7 \$3 \$4 \$4 sg13_lv_pmos W=4.0 L=0.13
.ENDS comp_5_split1

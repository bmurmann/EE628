* Extracted by KLayout with SG13G2 LVS runset on : 02/05/2024 06:37

* cell padring
* pin RES
* pin CK4
* pin CK5
* pin CK6
* pin IOVDD
* pin AVDD,IOVDD
* pin VDD
* pin res_c
* pin ck4_c
* pin ck5_c
* pin ck6_c
* pin IN6,PAD
* pin OUT6
* pin out6_c
* pin PADRES,in6_c
* pin IN5,PAD
* pin OUT5
* pin out5_c
* pin PADRES,in5_c
* pin IN4,PAD
* pin OUT4
* pin out4_c
* pin PADRES,in4_c
* pin PAD,VLO
* pin PADRES
* pin PAD,VHI
* pin PADRES
* pin IN3,PAD
* pin OUT3
* pin out3_c
* pin PADRES,in3_c
* pin IN2,PAD
* pin OUT2
* pin out2_c
* pin PADRES,in2_c
* pin IN1,PAD
* pin OUT1
* pin out1_c
* pin PADRES,in1_c
* pin PAD,VREF
* pin PADRES,vref_c
* pin PAD,VLDO
* pin ck3_c
* pin ck2_c
* pin ck1_c
* pin PADRES
* pin CK3
* pin CK2
* pin CK1
* pin IOVSS,VSS
.SUBCKT padring RES CK4 CK5 CK6 IOVDD AVDD|IOVDD VDD res_c ck4_c ck5_c ck6_c
+ IN6|PAD OUT6 out6_c PADRES|in6_c IN5|PAD OUT5 out5_c PADRES|in5_c IN4|PAD
+ OUT4 out4_c PADRES|in4_c PAD|VLO PADRES PAD|VHI PADRES$1 IN3|PAD OUT3 out3_c
+ PADRES|in3_c IN2|PAD OUT2 out2_c PADRES|in2_c IN1|PAD OUT1 out1_c
+ PADRES|in1_c PAD|VREF PADRES|vref_c PAD|VLDO ck3_c ck2_c ck1_c PADRES$2 CK3
+ CK2 CK1 IOVSS|VSS
* device instance $1 r0 *1 240.255,159.005 sg13_lv_nmos
M$1 res_c \$186 IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $2 r0 *1 440.255,159.005 sg13_lv_nmos
M$2 ck4_c \$187 IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $3 r0 *1 540.255,159.005 sg13_lv_nmos
M$3 ck5_c \$188 IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $4 r0 *1 640.255,159.005 sg13_lv_nmos
M$4 ck6_c \$189 IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $5 r0 *1 800.995,217.48 sg13_lv_nmos
M$5 \$237 out6_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $6 r0 *1 800.995,220.99 sg13_lv_nmos
M$6 \$264 out6_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $7 r0 *1 800.995,317.48 sg13_lv_nmos
M$7 \$350 out5_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $8 r0 *1 800.995,320.99 sg13_lv_nmos
M$8 \$377 out5_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $9 r0 *1 800.995,417.48 sg13_lv_nmos
M$9 \$463 out4_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $10 r0 *1 800.995,420.99 sg13_lv_nmos
M$10 \$490 out4_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $11 r0 *1 800.995,717.48 sg13_lv_nmos
M$11 \$776 out3_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $12 r0 *1 800.995,720.99 sg13_lv_nmos
M$12 \$803 out3_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $13 r0 *1 800.995,817.48 sg13_lv_nmos
M$13 \$889 out2_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $14 r0 *1 800.995,820.99 sg13_lv_nmos
M$14 \$916 out2_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $15 r0 *1 800.995,917.48 sg13_lv_nmos
M$15 \$1002 out1_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $16 r0 *1 800.995,920.99 sg13_lv_nmos
M$16 \$1029 out1_c IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $17 r0 *1 440.255,980.995 sg13_lv_nmos
M$17 ck3_c \$1092 IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $18 r0 *1 540.255,980.995 sg13_lv_nmos
M$18 ck2_c \$1093 IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $19 r0 *1 640.255,980.995 sg13_lv_nmos
M$19 ck1_c \$1094 IOVSS|VSS IOVSS|VSS sg13_lv_nmos W=2.7499999999999996
+ L=0.12999999999999995
* device instance $20 r0 *1 241.765,159.055 sg13_hv_nmos
M$20 IOVSS|VSS \$129 \$186 IOVSS|VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $21 r0 *1 441.765,159.055 sg13_hv_nmos
M$21 IOVSS|VSS \$130 \$187 IOVSS|VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $22 r0 *1 541.765,159.055 sg13_hv_nmos
M$22 IOVSS|VSS \$132 \$188 IOVSS|VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $23 r0 *1 641.765,159.055 sg13_hv_nmos
M$23 IOVSS|VSS \$133 \$189 IOVSS|VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $24 r0 *1 -169.05,205.52 sg13_hv_nmos
M$24 IOVSS|VSS \$227 IN6|PAD IOVSS|VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $44 r0 *1 949.05,214.58 sg13_hv_nmos
M$44 IOVSS|VSS \$253 OUT6 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $52 r0 *1 804.68,217.64 sg13_hv_nmos
M$52 \$238 out6_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $53 r0 *1 804.68,218.47 sg13_hv_nmos
M$53 IOVSS|VSS \$237 \$248 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $54 r0 *1 804.68,219.81 sg13_hv_nmos
M$54 IOVSS|VSS \$248 \$253 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $55 r0 *1 804.68,221.15 sg13_hv_nmos
M$55 \$265 out6_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $56 r0 *1 804.68,221.98 sg13_hv_nmos
M$56 IOVSS|VSS \$264 \$272 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $57 r0 *1 804.68,223.32 sg13_hv_nmos
M$57 IOVSS|VSS \$272 \$218 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $58 r0 *1 -169.05,305.52 sg13_hv_nmos
M$58 IOVSS|VSS \$340 IN5|PAD IOVSS|VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $78 r0 *1 949.05,314.58 sg13_hv_nmos
M$78 IOVSS|VSS \$366 OUT5 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $86 r0 *1 804.68,317.64 sg13_hv_nmos
M$86 \$351 out5_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $87 r0 *1 804.68,318.47 sg13_hv_nmos
M$87 IOVSS|VSS \$350 \$361 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $88 r0 *1 804.68,319.81 sg13_hv_nmos
M$88 IOVSS|VSS \$361 \$366 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $89 r0 *1 804.68,321.15 sg13_hv_nmos
M$89 \$378 out5_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $90 r0 *1 804.68,321.98 sg13_hv_nmos
M$90 IOVSS|VSS \$377 \$385 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $91 r0 *1 804.68,323.32 sg13_hv_nmos
M$91 IOVSS|VSS \$385 \$331 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $92 r0 *1 -169.05,405.52 sg13_hv_nmos
M$92 IOVSS|VSS \$453 IN4|PAD IOVSS|VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $112 r0 *1 949.05,414.58 sg13_hv_nmos
M$112 IOVSS|VSS \$479 OUT4 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $120 r0 *1 804.68,417.64 sg13_hv_nmos
M$120 \$464 out4_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $121 r0 *1 804.68,418.47 sg13_hv_nmos
M$121 IOVSS|VSS \$463 \$474 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $122 r0 *1 804.68,419.81 sg13_hv_nmos
M$122 IOVSS|VSS \$474 \$479 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $123 r0 *1 804.68,421.15 sg13_hv_nmos
M$123 \$491 out4_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $124 r0 *1 804.68,421.98 sg13_hv_nmos
M$124 IOVSS|VSS \$490 \$498 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $125 r0 *1 804.68,423.32 sg13_hv_nmos
M$125 IOVSS|VSS \$498 \$444 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $126 r0 *1 -169.05,505.52 sg13_hv_nmos
M$126 IOVSS|VSS \$568 PAD|VLO IOVSS|VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $146 r0 *1 879.21,583.22 sg13_hv_nmos
M$146 IOVSS|VSS \$627 \$626 IOVSS|VSS sg13_hv_nmos W=107.99999999999999
+ L=0.4999999999999999
* device instance $152 r0 *1 879.21,593 sg13_hv_nmos
M$152 IOVSS|VSS \$627 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=125.99999999999999
+ L=9.499999999999996
* device instance $172 r0 *1 934.53,588.155 sg13_hv_nmos
M$172 IOVSS|VSS \$626 IOVDD IOVSS|VSS sg13_hv_nmos W=756.7999999999977
+ L=0.5999999999999998
* device instance $344 r0 *1 -169.05,605.52 sg13_hv_nmos
M$344 IOVSS|VSS \$643 PAD|VHI IOVSS|VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $364 r0 *1 -169.05,705.52 sg13_hv_nmos
M$364 IOVSS|VSS \$766 IN3|PAD IOVSS|VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $384 r0 *1 949.05,714.58 sg13_hv_nmos
M$384 IOVSS|VSS \$792 OUT3 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $392 r0 *1 804.68,717.64 sg13_hv_nmos
M$392 \$777 out3_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $393 r0 *1 804.68,718.47 sg13_hv_nmos
M$393 IOVSS|VSS \$776 \$787 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $394 r0 *1 804.68,719.81 sg13_hv_nmos
M$394 IOVSS|VSS \$787 \$792 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $395 r0 *1 804.68,721.15 sg13_hv_nmos
M$395 \$804 out3_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $396 r0 *1 804.68,721.98 sg13_hv_nmos
M$396 IOVSS|VSS \$803 \$811 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $397 r0 *1 804.68,723.32 sg13_hv_nmos
M$397 IOVSS|VSS \$811 \$757 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $398 r0 *1 -169.05,805.52 sg13_hv_nmos
M$398 IOVSS|VSS \$879 IN2|PAD IOVSS|VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $418 r0 *1 949.05,814.58 sg13_hv_nmos
M$418 IOVSS|VSS \$905 OUT2 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $426 r0 *1 804.68,817.64 sg13_hv_nmos
M$426 \$890 out2_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $427 r0 *1 804.68,818.47 sg13_hv_nmos
M$427 IOVSS|VSS \$889 \$900 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $428 r0 *1 804.68,819.81 sg13_hv_nmos
M$428 IOVSS|VSS \$900 \$905 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $429 r0 *1 804.68,821.15 sg13_hv_nmos
M$429 \$917 out2_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $430 r0 *1 804.68,821.98 sg13_hv_nmos
M$430 IOVSS|VSS \$916 \$924 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $431 r0 *1 804.68,823.32 sg13_hv_nmos
M$431 IOVSS|VSS \$924 \$870 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $432 r0 *1 -169.05,905.52 sg13_hv_nmos
M$432 IOVSS|VSS \$992 IN1|PAD IOVSS|VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $452 r0 *1 949.05,914.58 sg13_hv_nmos
M$452 IOVSS|VSS \$1018 OUT1 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $460 r0 *1 804.68,917.64 sg13_hv_nmos
M$460 \$1003 out1_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $461 r0 *1 804.68,918.47 sg13_hv_nmos
M$461 IOVSS|VSS \$1002 \$1013 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $462 r0 *1 804.68,919.81 sg13_hv_nmos
M$462 IOVSS|VSS \$1013 \$1018 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $463 r0 *1 804.68,921.15 sg13_hv_nmos
M$463 \$1030 out1_c IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $464 r0 *1 804.68,921.98 sg13_hv_nmos
M$464 IOVSS|VSS \$1029 \$1037 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $465 r0 *1 804.68,923.32 sg13_hv_nmos
M$465 IOVSS|VSS \$1037 \$983 IOVSS|VSS sg13_hv_nmos W=1.8999999999999997
+ L=0.4499999999999999
* device instance $466 r0 *1 441.765,980.945 sg13_hv_nmos
M$466 IOVSS|VSS \$1095 \$1092 IOVSS|VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $467 r0 *1 541.765,980.945 sg13_hv_nmos
M$467 IOVSS|VSS \$1096 \$1093 IOVSS|VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $468 r0 *1 641.765,980.945 sg13_hv_nmos
M$468 IOVSS|VSS \$1097 \$1094 IOVSS|VSS sg13_hv_nmos W=2.6499999999999995
+ L=0.4499999999999999
* device instance $469 r0 *1 3.22,1059.21 sg13_hv_nmos
M$469 IOVSS|VSS \$1228 \$1169 IOVSS|VSS sg13_hv_nmos W=107.99999999999999
+ L=0.4999999999999999
* device instance $475 r0 *1 13,1059.21 sg13_hv_nmos
M$475 IOVSS|VSS \$1228 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=125.99999999999999
+ L=9.499999999999996
* device instance $482 r0 *1 303.22,1059.21 sg13_hv_nmos
M$482 IOVSS|VSS \$1229 \$1170 IOVSS|VSS sg13_hv_nmos W=107.99999999999999
+ L=0.4999999999999999
* device instance $488 r0 *1 313,1059.21 sg13_hv_nmos
M$488 IOVSS|VSS \$1229 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=125.99999999999999
+ L=9.499999999999996
* device instance $495 r0 *1 703.22,1059.21 sg13_hv_nmos
M$495 IOVSS|VSS \$1230 \$1171 IOVSS|VSS sg13_hv_nmos W=107.99999999999999
+ L=0.4999999999999999
* device instance $501 r0 *1 713,1059.21 sg13_hv_nmos
M$501 IOVSS|VSS \$1230 IOVSS|VSS IOVSS|VSS sg13_hv_nmos W=125.99999999999999
+ L=9.499999999999996
* device instance $547 r0 *1 8.155,1114.53 sg13_hv_nmos
M$547 IOVSS|VSS \$1169 \$1420 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $549 r0 *1 11.175,1114.53 sg13_hv_nmos
M$549 IOVSS|VSS \$1169 \$1421 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $551 r0 *1 14.195,1114.53 sg13_hv_nmos
M$551 IOVSS|VSS \$1169 \$1422 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $553 r0 *1 17.215,1114.53 sg13_hv_nmos
M$553 IOVSS|VSS \$1169 \$1423 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $555 r0 *1 20.235,1114.53 sg13_hv_nmos
M$555 IOVSS|VSS \$1169 \$1424 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $557 r0 *1 23.255,1114.53 sg13_hv_nmos
M$557 IOVSS|VSS \$1169 \$1425 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $559 r0 *1 26.275,1114.53 sg13_hv_nmos
M$559 IOVSS|VSS \$1169 \$1426 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $561 r0 *1 29.295,1114.53 sg13_hv_nmos
M$561 IOVSS|VSS \$1169 \$1427 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $563 r0 *1 32.315,1114.53 sg13_hv_nmos
M$563 IOVSS|VSS \$1169 \$1428 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $565 r0 *1 35.335,1114.53 sg13_hv_nmos
M$565 IOVSS|VSS \$1169 \$1429 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $567 r0 *1 38.355,1114.53 sg13_hv_nmos
M$567 IOVSS|VSS \$1169 \$1430 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $569 r0 *1 41.375,1114.53 sg13_hv_nmos
M$569 IOVSS|VSS \$1169 \$1431 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $571 r0 *1 44.395,1114.53 sg13_hv_nmos
M$571 IOVSS|VSS \$1169 \$1432 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $573 r0 *1 47.415,1114.53 sg13_hv_nmos
M$573 IOVSS|VSS \$1169 \$1433 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $575 r0 *1 50.435,1114.53 sg13_hv_nmos
M$575 IOVSS|VSS \$1169 \$1434 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $577 r0 *1 53.455,1114.53 sg13_hv_nmos
M$577 IOVSS|VSS \$1169 \$1435 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $579 r0 *1 56.475,1114.53 sg13_hv_nmos
M$579 IOVSS|VSS \$1169 \$1436 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $581 r0 *1 59.495,1114.53 sg13_hv_nmos
M$581 IOVSS|VSS \$1169 \$1437 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $583 r0 *1 62.515,1114.53 sg13_hv_nmos
M$583 IOVSS|VSS \$1169 \$1438 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $585 r0 *1 65.535,1114.53 sg13_hv_nmos
M$585 IOVSS|VSS \$1169 \$1439 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $587 r0 *1 68.555,1114.53 sg13_hv_nmos
M$587 IOVSS|VSS \$1169 \$1440 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $589 r0 *1 71.575,1114.53 sg13_hv_nmos
M$589 IOVSS|VSS \$1169 \$1441 IOVSS|VSS sg13_hv_nmos W=17.599999999999998
+ L=0.5999999999999998
* device instance $590 r0 *1 308.155,1114.53 sg13_hv_nmos
M$590 IOVSS|VSS \$1170 IOVDD IOVSS|VSS sg13_hv_nmos W=756.7999999999977
+ L=0.5999999999999998
* device instance $633 r0 *1 708.155,1114.53 sg13_hv_nmos
M$633 IOVSS|VSS \$1171 \$1442 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $635 r0 *1 711.175,1114.53 sg13_hv_nmos
M$635 IOVSS|VSS \$1171 \$1443 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $637 r0 *1 714.195,1114.53 sg13_hv_nmos
M$637 IOVSS|VSS \$1171 \$1444 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $639 r0 *1 717.215,1114.53 sg13_hv_nmos
M$639 IOVSS|VSS \$1171 \$1445 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $641 r0 *1 720.235,1114.53 sg13_hv_nmos
M$641 IOVSS|VSS \$1171 \$1446 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $643 r0 *1 723.255,1114.53 sg13_hv_nmos
M$643 IOVSS|VSS \$1171 \$1447 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $645 r0 *1 726.275,1114.53 sg13_hv_nmos
M$645 IOVSS|VSS \$1171 \$1448 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $647 r0 *1 729.295,1114.53 sg13_hv_nmos
M$647 IOVSS|VSS \$1171 \$1449 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $649 r0 *1 732.315,1114.53 sg13_hv_nmos
M$649 IOVSS|VSS \$1171 \$1450 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $651 r0 *1 735.335,1114.53 sg13_hv_nmos
M$651 IOVSS|VSS \$1171 \$1451 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $653 r0 *1 738.355,1114.53 sg13_hv_nmos
M$653 IOVSS|VSS \$1171 \$1452 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $655 r0 *1 741.375,1114.53 sg13_hv_nmos
M$655 IOVSS|VSS \$1171 \$1453 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $657 r0 *1 744.395,1114.53 sg13_hv_nmos
M$657 IOVSS|VSS \$1171 \$1454 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $659 r0 *1 747.415,1114.53 sg13_hv_nmos
M$659 IOVSS|VSS \$1171 \$1455 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $661 r0 *1 750.435,1114.53 sg13_hv_nmos
M$661 IOVSS|VSS \$1171 \$1456 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $663 r0 *1 753.455,1114.53 sg13_hv_nmos
M$663 IOVSS|VSS \$1171 \$1457 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $665 r0 *1 756.475,1114.53 sg13_hv_nmos
M$665 IOVSS|VSS \$1171 \$1458 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $667 r0 *1 759.495,1114.53 sg13_hv_nmos
M$667 IOVSS|VSS \$1171 \$1459 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $669 r0 *1 762.515,1114.53 sg13_hv_nmos
M$669 IOVSS|VSS \$1171 \$1460 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $671 r0 *1 765.535,1114.53 sg13_hv_nmos
M$671 IOVSS|VSS \$1171 \$1461 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $673 r0 *1 768.555,1114.53 sg13_hv_nmos
M$673 IOVSS|VSS \$1171 \$1462 IOVSS|VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999998
* device instance $675 r0 *1 771.575,1114.53 sg13_hv_nmos
M$675 IOVSS|VSS \$1171 \$1463 IOVSS|VSS sg13_hv_nmos W=17.599999999999998
+ L=0.5999999999999998
* device instance $977 r0 *1 125.52,1129.05 sg13_hv_nmos
M$977 IOVSS|VSS \$1501 PAD|VREF IOVSS|VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $997 r0 *1 225.52,1129.05 sg13_hv_nmos
M$997 IOVSS|VSS \$1502 PAD|VLDO IOVSS|VSS sg13_hv_nmos W=88.00000000000001
+ L=0.5999999999999998
* device instance $1103 r0 *1 240.255,163.995 sg13_lv_pmos
M$1103 res_c \$186 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1104 r0 *1 440.255,163.995 sg13_lv_pmos
M$1104 ck4_c \$187 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1105 r0 *1 540.255,163.995 sg13_lv_pmos
M$1105 ck5_c \$188 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1106 r0 *1 640.255,163.995 sg13_lv_pmos
M$1106 ck6_c \$189 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1107 r0 *1 796.005,217.48 sg13_lv_pmos
M$1107 \$237 out6_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1108 r0 *1 796.005,220.99 sg13_lv_pmos
M$1108 \$264 out6_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1109 r0 *1 796.005,317.48 sg13_lv_pmos
M$1109 \$350 out5_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1110 r0 *1 796.005,320.99 sg13_lv_pmos
M$1110 \$377 out5_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1111 r0 *1 796.005,417.48 sg13_lv_pmos
M$1111 \$463 out4_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1112 r0 *1 796.005,420.99 sg13_lv_pmos
M$1112 \$490 out4_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1113 r0 *1 796.005,717.48 sg13_lv_pmos
M$1113 \$776 out3_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1114 r0 *1 796.005,720.99 sg13_lv_pmos
M$1114 \$803 out3_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1115 r0 *1 796.005,817.48 sg13_lv_pmos
M$1115 \$889 out2_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1116 r0 *1 796.005,820.99 sg13_lv_pmos
M$1116 \$916 out2_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1117 r0 *1 796.005,917.48 sg13_lv_pmos
M$1117 \$1002 out1_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1118 r0 *1 796.005,920.99 sg13_lv_pmos
M$1118 \$1029 out1_c VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1119 r0 *1 440.255,976.005 sg13_lv_pmos
M$1119 ck3_c \$1092 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1120 r0 *1 540.255,976.005 sg13_lv_pmos
M$1120 ck2_c \$1093 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1121 r0 *1 640.255,976.005 sg13_lv_pmos
M$1121 ck1_c \$1094 VDD VDD sg13_lv_pmos W=4.749999999999999
+ L=0.12999999999999998
* device instance $1122 r0 *1 241.765,163.945 sg13_hv_pmos
M$1122 VDD \$129 \$186 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1123 r0 *1 441.765,163.945 sg13_hv_pmos
M$1123 VDD \$130 \$187 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1124 r0 *1 541.765,163.945 sg13_hv_pmos
M$1124 VDD \$132 \$188 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1125 r0 *1 641.765,163.945 sg13_hv_pmos
M$1125 VDD \$133 \$189 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1126 r0 *1 -108.92,205.52 sg13_hv_pmos
M$1126 AVDD|IOVDD \$228 IN6|PAD AVDD|IOVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1166 r0 *1 881.82,214.58 sg13_hv_pmos
M$1166 IOVDD \$218 OUT6 IOVDD sg13_hv_pmos W=106.55999999999996
+ L=0.5999999999999999
* device instance $1182 r0 *1 808.82,217.64 sg13_hv_pmos
M$1182 \$238 \$248 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1183 r0 *1 808.82,218.47 sg13_hv_pmos
M$1183 IOVDD \$238 \$248 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1184 r0 *1 808.82,219.81 sg13_hv_pmos
M$1184 IOVDD \$248 \$253 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1185 r0 *1 808.82,221.15 sg13_hv_pmos
M$1185 \$265 \$272 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1186 r0 *1 808.82,221.98 sg13_hv_pmos
M$1186 IOVDD \$265 \$272 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1187 r0 *1 808.82,223.32 sg13_hv_pmos
M$1187 IOVDD \$272 \$218 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1188 r0 *1 -108.92,305.52 sg13_hv_pmos
M$1188 AVDD|IOVDD \$341 IN5|PAD AVDD|IOVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1228 r0 *1 881.82,314.58 sg13_hv_pmos
M$1228 IOVDD \$331 OUT5 IOVDD sg13_hv_pmos W=106.55999999999996
+ L=0.5999999999999999
* device instance $1244 r0 *1 808.82,317.64 sg13_hv_pmos
M$1244 \$351 \$361 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1245 r0 *1 808.82,318.47 sg13_hv_pmos
M$1245 IOVDD \$351 \$361 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1246 r0 *1 808.82,319.81 sg13_hv_pmos
M$1246 IOVDD \$361 \$366 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1247 r0 *1 808.82,321.15 sg13_hv_pmos
M$1247 \$378 \$385 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1248 r0 *1 808.82,321.98 sg13_hv_pmos
M$1248 IOVDD \$378 \$385 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1249 r0 *1 808.82,323.32 sg13_hv_pmos
M$1249 IOVDD \$385 \$331 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1250 r0 *1 -108.92,405.52 sg13_hv_pmos
M$1250 AVDD|IOVDD \$454 IN4|PAD AVDD|IOVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1290 r0 *1 881.82,414.58 sg13_hv_pmos
M$1290 IOVDD \$444 OUT4 IOVDD sg13_hv_pmos W=106.55999999999996
+ L=0.5999999999999999
* device instance $1306 r0 *1 808.82,417.64 sg13_hv_pmos
M$1306 \$464 \$474 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1307 r0 *1 808.82,418.47 sg13_hv_pmos
M$1307 IOVDD \$464 \$474 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1308 r0 *1 808.82,419.81 sg13_hv_pmos
M$1308 IOVDD \$474 \$479 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1309 r0 *1 808.82,421.15 sg13_hv_pmos
M$1309 \$491 \$498 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1310 r0 *1 808.82,421.98 sg13_hv_pmos
M$1310 IOVDD \$491 \$498 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1311 r0 *1 808.82,423.32 sg13_hv_pmos
M$1311 IOVDD \$498 \$444 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1312 r0 *1 -108.92,505.52 sg13_hv_pmos
M$1312 AVDD|IOVDD \$569 PAD|VLO AVDD|IOVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1352 r0 *1 865.09,598.44 sg13_hv_pmos
M$1352 IOVDD \$627 \$626 IOVDD sg13_hv_pmos W=349.99999999999994
+ L=0.4999999999999999
* device instance $1402 r0 *1 -108.92,605.52 sg13_hv_pmos
M$1402 AVDD|IOVDD \$644 PAD|VHI AVDD|IOVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1442 r0 *1 -108.92,705.52 sg13_hv_pmos
M$1442 AVDD|IOVDD \$767 IN3|PAD AVDD|IOVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1482 r0 *1 881.82,714.58 sg13_hv_pmos
M$1482 IOVDD \$757 OUT3 IOVDD sg13_hv_pmos W=106.55999999999996
+ L=0.5999999999999999
* device instance $1498 r0 *1 808.82,717.64 sg13_hv_pmos
M$1498 \$777 \$787 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1499 r0 *1 808.82,718.47 sg13_hv_pmos
M$1499 IOVDD \$777 \$787 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1500 r0 *1 808.82,719.81 sg13_hv_pmos
M$1500 IOVDD \$787 \$792 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1501 r0 *1 808.82,721.15 sg13_hv_pmos
M$1501 \$804 \$811 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1502 r0 *1 808.82,721.98 sg13_hv_pmos
M$1502 IOVDD \$804 \$811 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1503 r0 *1 808.82,723.32 sg13_hv_pmos
M$1503 IOVDD \$811 \$757 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1504 r0 *1 -108.92,805.52 sg13_hv_pmos
M$1504 AVDD|IOVDD \$880 IN2|PAD AVDD|IOVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1544 r0 *1 881.82,814.58 sg13_hv_pmos
M$1544 IOVDD \$870 OUT2 IOVDD sg13_hv_pmos W=106.55999999999996
+ L=0.5999999999999999
* device instance $1560 r0 *1 808.82,817.64 sg13_hv_pmos
M$1560 \$890 \$900 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1561 r0 *1 808.82,818.47 sg13_hv_pmos
M$1561 IOVDD \$890 \$900 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1562 r0 *1 808.82,819.81 sg13_hv_pmos
M$1562 IOVDD \$900 \$905 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1563 r0 *1 808.82,821.15 sg13_hv_pmos
M$1563 \$917 \$924 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1564 r0 *1 808.82,821.98 sg13_hv_pmos
M$1564 IOVDD \$917 \$924 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1565 r0 *1 808.82,823.32 sg13_hv_pmos
M$1565 IOVDD \$924 \$870 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1566 r0 *1 -108.92,905.52 sg13_hv_pmos
M$1566 AVDD|IOVDD \$993 IN1|PAD AVDD|IOVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1606 r0 *1 881.82,914.58 sg13_hv_pmos
M$1606 IOVDD \$983 OUT1 IOVDD sg13_hv_pmos W=106.55999999999996
+ L=0.5999999999999999
* device instance $1622 r0 *1 808.82,917.64 sg13_hv_pmos
M$1622 \$1003 \$1013 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1623 r0 *1 808.82,918.47 sg13_hv_pmos
M$1623 IOVDD \$1003 \$1013 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1624 r0 *1 808.82,919.81 sg13_hv_pmos
M$1624 IOVDD \$1013 \$1018 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1625 r0 *1 808.82,921.15 sg13_hv_pmos
M$1625 \$1030 \$1037 IOVDD IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1626 r0 *1 808.82,921.98 sg13_hv_pmos
M$1626 IOVDD \$1030 \$1037 IOVDD sg13_hv_pmos W=0.29999999999999993
+ L=0.44999999999999984
* device instance $1627 r0 *1 808.82,923.32 sg13_hv_pmos
M$1627 IOVDD \$1037 \$983 IOVDD sg13_hv_pmos W=3.899999999999999
+ L=0.4499999999999999
* device instance $1628 r0 *1 441.765,976.055 sg13_hv_pmos
M$1628 VDD \$1095 \$1092 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1629 r0 *1 541.765,976.055 sg13_hv_pmos
M$1629 VDD \$1096 \$1093 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1630 r0 *1 641.765,976.055 sg13_hv_pmos
M$1630 VDD \$1097 \$1094 VDD sg13_hv_pmos W=4.6499999999999995
+ L=0.44999999999999984
* device instance $1631 r0 *1 18.44,1045.09 sg13_hv_pmos
M$1631 AVDD|IOVDD \$1228 \$1169 AVDD|IOVDD sg13_hv_pmos W=349.99999999999994
+ L=0.4999999999999999
* device instance $1681 r0 *1 318.44,1045.09 sg13_hv_pmos
M$1681 IOVDD \$1229 \$1170 IOVDD sg13_hv_pmos W=349.99999999999994
+ L=0.4999999999999999
* device instance $1731 r0 *1 718.44,1045.09 sg13_hv_pmos
M$1731 IOVDD \$1230 \$1171 IOVDD sg13_hv_pmos W=349.99999999999994
+ L=0.4999999999999999
* device instance $1781 r0 *1 125.52,1061.82 sg13_hv_pmos
M$1781 AVDD|IOVDD \$1186 PAD|VREF AVDD|IOVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1821 r0 *1 225.52,1061.82 sg13_hv_pmos
M$1821 AVDD|IOVDD \$1187 PAD|VLDO AVDD|IOVDD sg13_hv_pmos W=266.3999999999999
+ L=0.5999999999999999
* device instance $1861 r0 *1 4.54,24.19 dantenna
D$1861 IOVSS|VSS IOVSS|VSS dantenna A=35.0028 P=58.08 m=10
* device instance $1865 r0 *1 204.54,24.19 dantenna
D$1865 IOVSS|VSS RES dantenna A=35.0028 P=58.08 m=2
* device instance $1869 r0 *1 404.54,24.19 dantenna
D$1869 IOVSS|VSS CK4 dantenna A=35.0028 P=58.08 m=2
* device instance $1871 r0 *1 504.54,24.19 dantenna
D$1871 IOVSS|VSS CK5 dantenna A=35.0028 P=58.08 m=2
* device instance $1873 r0 *1 604.54,24.19 dantenna
D$1873 IOVSS|VSS CK6 dantenna A=35.0028 P=58.08 m=2
* device instance $1877 r0 *1 -159.56,320 dantenna
D$1877 IOVSS|VSS IN5|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1878 r0 *1 -159.56,220 dantenna
D$1878 IOVSS|VSS IN6|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1881 r0 *1 -37.46,337.63 dantenna
D$1881 IOVSS|VSS PADRES|in5_c dantenna A=1.984 P=7.48 m=1
* device instance $1882 r0 *1 -37.46,237.63 dantenna
D$1882 IOVSS|VSS PADRES|in6_c dantenna A=1.984 P=7.48 m=1
* device instance $1883 r0 *1 245.225,142.54 dantenna
D$1883 IOVSS|VSS \$129 dantenna A=1.984 P=7.48 m=1
* device instance $1884 r0 *1 445.225,142.54 dantenna
D$1884 IOVSS|VSS \$130 dantenna A=1.984 P=7.48 m=1
* device instance $1885 r0 *1 545.225,142.54 dantenna
D$1885 IOVSS|VSS \$132 dantenna A=1.984 P=7.48 m=1
* device instance $1886 r0 *1 645.225,142.54 dantenna
D$1886 IOVSS|VSS \$133 dantenna A=1.984 P=7.48 m=1
* device instance $1887 r0 *1 935.06,220 dantenna
D$1887 IOVSS|VSS OUT6 dantenna A=35.0028 P=58.08 m=2
* device instance $1888 r0 *1 935.06,320 dantenna
D$1888 IOVSS|VSS OUT5 dantenna A=35.0028 P=58.08 m=2
* device instance $1891 r0 *1 947.17,297.975 dantenna
D$1891 IOVSS|VSS \$366 dantenna A=0.192 P=1.88 m=1
* device instance $1892 r0 *1 947.17,197.975 dantenna
D$1892 IOVSS|VSS \$253 dantenna A=0.192 P=1.88 m=1
* device instance $1893 r0 *1 947.17,397.975 dantenna
D$1893 IOVSS|VSS \$479 dantenna A=0.192 P=1.88 m=1
* device instance $1894 r0 *1 -159.56,420 dantenna
D$1894 IOVSS|VSS IN4|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1896 r0 *1 935.06,420 dantenna
D$1896 IOVSS|VSS OUT4 dantenna A=35.0028 P=58.08 m=2
* device instance $1898 r0 *1 -37.46,437.63 dantenna
D$1898 IOVSS|VSS PADRES|in4_c dantenna A=1.984 P=7.48 m=1
* device instance $1901 r0 *1 -159.56,520 dantenna
D$1901 IOVSS|VSS PAD|VLO dantenna A=35.0028 P=58.08 m=2
* device instance $1903 r0 *1 -37.46,537.63 dantenna
D$1903 IOVSS|VSS PADRES dantenna A=1.984 P=7.48 m=1
* device instance $1904 r0 *1 932.65,584.765 dantenna
D$1904 IOVSS|VSS \$626 dantenna A=0.192 P=1.88 m=1
* device instance $1905 r0 *1 -159.56,620 dantenna
D$1905 IOVSS|VSS PAD|VHI dantenna A=35.0028 P=58.08 m=2
* device instance $1907 r0 *1 -37.46,637.63 dantenna
D$1907 IOVSS|VSS PADRES$1 dantenna A=1.984 P=7.48 m=1
* device instance $1908 r0 *1 947.17,697.975 dantenna
D$1908 IOVSS|VSS \$792 dantenna A=0.192 P=1.88 m=1
* device instance $1909 r0 *1 -159.56,720 dantenna
D$1909 IOVSS|VSS IN3|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1911 r0 *1 935.06,720 dantenna
D$1911 IOVSS|VSS OUT3 dantenna A=35.0028 P=58.08 m=2
* device instance $1913 r0 *1 -37.46,737.63 dantenna
D$1913 IOVSS|VSS PADRES|in3_c dantenna A=1.984 P=7.48 m=1
* device instance $1914 r0 *1 947.17,797.975 dantenna
D$1914 IOVSS|VSS \$905 dantenna A=0.192 P=1.88 m=1
* device instance $1915 r0 *1 -159.56,820 dantenna
D$1915 IOVSS|VSS IN2|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1917 r0 *1 935.06,820 dantenna
D$1917 IOVSS|VSS OUT2 dantenna A=35.0028 P=58.08 m=2
* device instance $1919 r0 *1 -37.46,837.63 dantenna
D$1919 IOVSS|VSS PADRES|in2_c dantenna A=1.984 P=7.48 m=1
* device instance $1920 r0 *1 947.17,897.975 dantenna
D$1920 IOVSS|VSS \$1018 dantenna A=0.192 P=1.88 m=1
* device instance $1921 r0 *1 -159.56,920 dantenna
D$1921 IOVSS|VSS IN1|PAD dantenna A=35.0028 P=58.08 m=2
* device instance $1923 r0 *1 935.06,920 dantenna
D$1923 IOVSS|VSS OUT1 dantenna A=35.0028 P=58.08 m=2
* device instance $1925 r0 *1 -37.46,937.63 dantenna
D$1925 IOVSS|VSS PADRES|in1_c dantenna A=1.984 P=7.48 m=1
* device instance $1926 r0 *1 157.63,997.46 dantenna
D$1926 IOVSS|VSS PADRES|vref_c dantenna A=1.984 P=7.48 m=1
* device instance $1927 r0 *1 257.63,997.46 dantenna
D$1927 IOVSS|VSS PADRES$2 dantenna A=1.984 P=7.48 m=1
* device instance $1928 r0 *1 445.225,997.46 dantenna
D$1928 IOVSS|VSS \$1095 dantenna A=1.984 P=7.48 m=1
* device instance $1929 r0 *1 545.225,997.46 dantenna
D$1929 IOVSS|VSS \$1096 dantenna A=1.984 P=7.48 m=1
* device instance $1930 r0 *1 645.225,997.46 dantenna
D$1930 IOVSS|VSS \$1097 dantenna A=1.984 P=7.48 m=1
* device instance $1931 r0 *1 404.54,1115.81 dantenna
D$1931 IOVSS|VSS CK3 dantenna A=35.0028 P=58.08 m=2
* device instance $1933 r0 *1 504.54,1115.81 dantenna
D$1933 IOVSS|VSS CK2 dantenna A=35.0028 P=58.08 m=2
* device instance $1935 r0 *1 604.54,1115.81 dantenna
D$1935 IOVSS|VSS CK1 dantenna A=35.0028 P=58.08 m=2
* device instance $1937 r0 *1 4.765,1112.65 dantenna
D$1937 IOVSS|VSS \$1169 dantenna A=0.192 P=1.88 m=1
* device instance $1938 r0 *1 140,1115.06 dantenna
D$1938 IOVSS|VSS PAD|VREF dantenna A=35.0028 P=58.08 m=2
* device instance $1939 r0 *1 240,1115.06 dantenna
D$1939 IOVSS|VSS PAD|VLDO dantenna A=35.0028 P=58.08 m=2
* device instance $1940 r0 *1 304.765,1112.65 dantenna
D$1940 IOVSS|VSS \$1170 dantenna A=0.192 P=1.88 m=1
* device instance $1941 r0 *1 704.765,1112.65 dantenna
D$1941 IOVSS|VSS \$1171 dantenna A=0.192 P=1.88 m=1
* device instance $1944 r0 *1 4.54,83.19 dpantenna
D$1944 IOVSS|VSS AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=4
* device instance $1948 r0 *1 204.54,83.19 dpantenna
D$1948 RES IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1950 r0 *1 304.54,83.19 dpantenna
D$1950 IOVSS|VSS IOVDD dpantenna A=35.0028 P=58.08 m=6
* device instance $1952 r0 *1 404.54,83.19 dpantenna
D$1952 CK4 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1954 r0 *1 504.54,83.19 dpantenna
D$1954 CK5 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1956 r0 *1 604.54,83.19 dpantenna
D$1956 CK6 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1960 r0 *1 -124.04,320 dpantenna
D$1960 IN5|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1961 r0 *1 -124.04,220 dpantenna
D$1961 IN6|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1964 r0 *1 -32.49,335.46 dpantenna
D$1964 PADRES|in5_c AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1965 r0 *1 -32.49,235.46 dpantenna
D$1965 PADRES|in6_c AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1966 r0 *1 243.055,147.51 dpantenna
D$1966 \$129 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1967 r0 *1 443.055,147.51 dpantenna
D$1967 \$130 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1968 r0 *1 543.055,147.51 dpantenna
D$1968 \$132 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1969 r0 *1 643.055,147.51 dpantenna
D$1969 \$133 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1970 r0 *1 878.81,197.975 dpantenna
D$1970 \$218 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $1971 r0 *1 878.81,297.975 dpantenna
D$1971 \$331 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $1972 r0 *1 899.54,320 dpantenna
D$1972 OUT5 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1973 r0 *1 899.54,220 dpantenna
D$1973 OUT6 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1976 r0 *1 -124.04,420 dpantenna
D$1976 IN4|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1978 r0 *1 878.81,397.975 dpantenna
D$1978 \$444 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $1979 r0 *1 899.54,420 dpantenna
D$1979 OUT4 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1981 r0 *1 -32.49,435.46 dpantenna
D$1981 PADRES|in4_c AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1984 r0 *1 -124.04,520 dpantenna
D$1984 PAD|VLO AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1986 r0 *1 -32.49,535.46 dpantenna
D$1986 PADRES AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1987 r0 *1 -124.04,620 dpantenna
D$1987 PAD|VHI AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1989 r0 *1 -32.49,635.46 dpantenna
D$1989 PADRES$1 AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1990 r0 *1 878.81,697.975 dpantenna
D$1990 \$757 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $1991 r0 *1 -124.04,720 dpantenna
D$1991 IN3|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1993 r0 *1 899.54,720 dpantenna
D$1993 OUT3 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1995 r0 *1 -32.49,735.46 dpantenna
D$1995 PADRES|in3_c AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $1996 r0 *1 878.81,797.975 dpantenna
D$1996 \$870 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $1997 r0 *1 -124.04,820 dpantenna
D$1997 IN2|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $1999 r0 *1 899.54,820 dpantenna
D$1999 OUT2 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2001 r0 *1 -32.49,835.46 dpantenna
D$2001 PADRES|in2_c AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2002 r0 *1 878.81,897.975 dpantenna
D$2002 \$983 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $2003 r0 *1 -124.04,920 dpantenna
D$2003 IN1|PAD AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2005 r0 *1 899.54,920 dpantenna
D$2005 OUT1 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2007 r0 *1 -32.49,935.46 dpantenna
D$2007 PADRES|in1_c AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2008 r0 *1 155.46,992.49 dpantenna
D$2008 PADRES|vref_c AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2009 r0 *1 255.46,992.49 dpantenna
D$2009 PADRES$2 AVDD|IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2010 r0 *1 443.055,992.49 dpantenna
D$2010 \$1095 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2011 r0 *1 543.055,992.49 dpantenna
D$2011 \$1096 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2012 r0 *1 643.055,992.49 dpantenna
D$2012 \$1097 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $2013 r0 *1 404.54,1056.81 dpantenna
D$2013 CK3 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2015 r0 *1 504.54,1056.81 dpantenna
D$2015 CK2 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2017 r0 *1 604.54,1056.81 dpantenna
D$2017 CK1 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2019 r0 *1 140,1084.04 dpantenna
D$2019 PAD|VREF AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2021 r0 *1 240,1084.04 dpantenna
D$2021 PAD|VLDO AVDD|IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $2023 r0 *1 240.685,141.11 res_rppd
R$2023 RES \$129 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $2024 r0 *1 440.685,141.11 res_rppd
R$2024 CK4 \$130 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $2025 r0 *1 540.685,141.11 res_rppd
R$2025 CK5 \$132 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $2026 r0 *1 640.685,141.11 res_rppd
R$2026 CK6 \$133 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $2027 r0 *1 -171.25,246.305 res_rppd
R$2027 IOVSS|VSS \$227 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2028 r0 *1 -112.25,246.305 res_rppd
R$2028 AVDD|IOVDD \$228 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $2029 r0 *1 -38.89,233.09 res_rppd
R$2029 IN6|PAD PADRES|in6_c res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $2030 r0 *1 -171.25,346.305 res_rppd
R$2030 IOVSS|VSS \$340 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2031 r0 *1 -112.25,346.305 res_rppd
R$2031 AVDD|IOVDD \$341 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $2032 r0 *1 -38.89,333.09 res_rppd
R$2032 IN5|PAD PADRES|in5_c res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $2033 r0 *1 -171.25,446.305 res_rppd
R$2033 IOVSS|VSS \$453 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2034 r0 *1 -112.25,446.305 res_rppd
R$2034 AVDD|IOVDD \$454 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $2035 r0 *1 -38.89,433.09 res_rppd
R$2035 IN4|PAD PADRES|in4_c res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $2036 r0 *1 -171.25,546.305 res_rppd
R$2036 IOVSS|VSS \$568 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2037 r0 *1 -112.25,546.305 res_rppd
R$2037 AVDD|IOVDD \$569 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $2038 r0 *1 -38.89,533.09 res_rppd
R$2038 PAD|VLO PADRES res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $2040 r0 *1 901.86,600.525 res_rppd
R$2040 \$635 \$633 res_rppd w=0.9999999999999998 l=79.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2043 r0 *1 901.86,605.475 res_rppd
R$2043 \$640 \$645 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2046 r0 *1 901.86,610.425 res_rppd
R$2046 \$655 \$651 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2048 r0 *1 901.86,613.725 res_rppd
R$2048 \$661 \$657 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2050 r0 *1 901.86,617.025 res_rppd
R$2050 \$667 \$663 res_rppd w=0.9999999999999998 l=79.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2053 r0 *1 901.86,621.975 res_rppd
R$2053 \$675 \$683 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2055 r0 *1 901.86,625.275 res_rppd
R$2055 \$685 \$689 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2057 r0 *1 901.86,628.575 res_rppd
R$2057 \$691 \$695 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2059 r0 *1 901.86,631.875 res_rppd
R$2059 \$697 \$701 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2060 r0 *1 -38.89,633.09 res_rppd
R$2060 PAD|VHI PADRES$1 res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $2063 r0 *1 901.86,636.825 res_rppd
R$2063 \$726 \$715 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2065 r0 *1 901.86,640.125 res_rppd
R$2065 \$627 \$731 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2066 r0 *1 -171.25,646.305 res_rppd
R$2066 IOVSS|VSS \$643 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2067 r0 *1 -112.25,646.305 res_rppd
R$2067 AVDD|IOVDD \$644 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $2068 r0 *1 -171.25,746.305 res_rppd
R$2068 IOVSS|VSS \$766 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2069 r0 *1 -112.25,746.305 res_rppd
R$2069 AVDD|IOVDD \$767 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $2070 r0 *1 -38.89,733.09 res_rppd
R$2070 IN3|PAD PADRES|in3_c res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $2071 r0 *1 -171.25,846.305 res_rppd
R$2071 IOVSS|VSS \$879 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2072 r0 *1 -112.25,846.305 res_rppd
R$2072 AVDD|IOVDD \$880 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $2073 r0 *1 -38.89,833.09 res_rppd
R$2073 IN2|PAD PADRES|in2_c res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $2074 r0 *1 -171.25,946.305 res_rppd
R$2074 IOVSS|VSS \$992 res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2075 r0 *1 -112.25,946.305 res_rppd
R$2075 AVDD|IOVDD \$993 res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $2076 r0 *1 -38.89,933.09 res_rppd
R$2076 IN1|PAD PADRES|in1_c res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $2077 r0 *1 153.09,996.03 res_rppd
R$2077 PADRES|vref_c PAD|VREF res_rppd w=0.9999999999999998
+ l=1.9999999999999996 b=0.0 ps=0.0 m=1.0
* device instance $2078 r0 *1 253.09,996.03 res_rppd
R$2078 PADRES$2 PAD|VLDO res_rppd w=0.9999999999999998 l=1.9999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $2079 r0 *1 440.685,996.03 res_rppd
R$2079 \$1095 CK3 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $2080 r0 *1 540.685,996.03 res_rppd
R$2080 \$1096 CK2 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $2081 r0 *1 640.685,996.03 res_rppd
R$2081 \$1097 CK1 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $2082 r0 *1 166.305,1058.49 res_rppd
R$2082 \$1186 AVDD|IOVDD res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $2083 r0 *1 266.305,1058.49 res_rppd
R$2083 \$1187 AVDD|IOVDD res_rppd w=0.4999999999999999 l=12.899999999999997
+ b=0.0 ps=0.0 m=1.0
* device instance $2084 r0 *1 18.875,1081.86 res_rppd
R$2084 AVDD|IOVDD \$1378 res_rppd w=0.9999999999999998 l=19.999999999999996
+ b=0.0 ps=0.0 m=1.0
* device instance $2085 r0 *1 20.525,1081.86 res_rppd
R$2085 \$1253 \$1378 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2087 r0 *1 23.825,1081.86 res_rppd
R$2087 \$1254 \$1379 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2089 r0 *1 27.125,1081.86 res_rppd
R$2089 \$1255 \$1380 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2091 r0 *1 30.425,1081.86 res_rppd
R$2091 \$1256 \$1381 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2093 r0 *1 33.725,1081.86 res_rppd
R$2093 \$1257 \$1382 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2097 r0 *1 40.325,1081.86 res_rppd
R$2097 \$1259 \$1384 res_rppd w=0.9999999999999998 l=79.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2100 r0 *1 45.275,1081.86 res_rppd
R$2100 \$1260 \$1386 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2103 r0 *1 50.225,1081.86 res_rppd
R$2103 \$1262 \$1387 res_rppd w=0.9999999999999998 l=79.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2105 r0 *1 53.525,1081.86 res_rppd
R$2105 \$1263 \$1388 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2107 r0 *1 56.825,1081.86 res_rppd
R$2107 \$1264 \$1389 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2109 r0 *1 60.125,1081.86 res_rppd
R$2109 \$1228 \$1390 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $2110 r0 *1 318.875,1081.86 res_rppd
R$2110 IOVDD \$1391 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $2111 r0 *1 320.525,1081.86 res_rppd
R$2111 \$1265 \$1391 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2113 r0 *1 323.825,1081.86 res_rppd
R$2113 \$1266 \$1392 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2115 r0 *1 327.125,1081.86 res_rppd
R$2115 \$1267 \$1393 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2117 r0 *1 330.425,1081.86 res_rppd
R$2117 \$1268 \$1394 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2120 r0 *1 335.375,1081.86 res_rppd
R$2120 \$1269 \$1396 res_rppd w=0.9999999999999998 l=79.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2123 r0 *1 340.325,1081.86 res_rppd
R$2123 \$1271 \$1397 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2125 r0 *1 343.625,1081.86 res_rppd
R$2125 \$1272 \$1398 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2127 r0 *1 346.925,1081.86 res_rppd
R$2127 \$1273 \$1399 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2131 r0 *1 353.525,1081.86 res_rppd
R$2131 \$1275 \$1401 res_rppd w=0.9999999999999998 l=79.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2133 r0 *1 356.825,1081.86 res_rppd
R$2133 \$1276 \$1402 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2135 r0 *1 360.125,1081.86 res_rppd
R$2135 \$1229 \$1403 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $2136 r0 *1 718.875,1081.86 res_rppd
R$2136 VDD \$1404 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $2139 r0 *1 723.825,1081.86 res_rppd
R$2139 \$1278 \$1405 res_rppd w=0.9999999999999998 l=79.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2142 r0 *1 728.775,1081.86 res_rppd
R$2142 \$1279 \$1407 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2144 r0 *1 732.075,1081.86 res_rppd
R$2144 \$1280 \$1408 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2146 r0 *1 735.375,1081.86 res_rppd
R$2146 \$1281 \$1409 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2148 r0 *1 738.675,1081.86 res_rppd
R$2148 \$1282 \$1410 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2150 r0 *1 741.975,1081.86 res_rppd
R$2150 \$1283 \$1411 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2152 r0 *1 745.275,1081.86 res_rppd
R$2152 \$1284 \$1412 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2155 r0 *1 750.225,1081.86 res_rppd
R$2155 \$1286 \$1413 res_rppd w=0.9999999999999998 l=79.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2158 r0 *1 755.175,1081.86 res_rppd
R$2158 \$1287 \$1415 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2160 r0 *1 758.475,1081.86 res_rppd
R$2160 \$1288 \$1416 res_rppd w=0.9999999999999998 l=39.99999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2161 r0 *1 760.125,1081.86 res_rppd
R$2161 \$1230 \$1416 res_rppd w=0.9999999999999998 l=19.999999999999996 b=0.0
+ ps=0.0 m=1.0
* device instance $2162 r0 *1 166.305,1126.85 res_rppd
R$2162 \$1501 IOVSS|VSS res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
* device instance $2163 r0 *1 266.305,1126.85 res_rppd
R$2163 \$1502 IOVSS|VSS res_rppd w=0.4999999999999999 l=3.539999999999999 b=0.0
+ ps=0.0 m=1.0
.ENDS padring

* Extracted by KLayout with SG13G2 LVS runset on : 03/05/2024 03:00

* cell sg13g2_SecondaryProtection
.SUBCKT sg13g2_SecondaryProtection
* device instance $1 r0 *1 5.48,2.37 dantenna
D$1 sub!$2 CORE dantenna A=1.984 P=7.48 m=1
* device instance $2 r0 *1 3.31,7.34 dpantenna
D$2 CORE \$10 dpantenna A=3.1872 P=11.24 m=1
* device instance $3 r0 *1 0.94,0.94 rppd
R$3 PAD CORE rppd w=1 l=2 ps=0 b=0 m=1
.ENDS sg13g2_SecondaryProtection

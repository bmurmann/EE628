* Extracted by KLayout with SG13G2 LVS runset on : 04/05/2024 17:50

* cell lvs_test
* pin vout
* pin vdda
* pin vss
.SUBCKT lvs_test vout vdda vss
* device instance $1 r0 *1 5.68,8.49 sg13_lv_nmos
M$1 vss \$4 \$1 vss sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $2 r0 *1 13.023,16.328 sg13_lv_nmos
M$2 vss \$1 vout vss sg13_lv_nmos W=0.9999999999999998 L=0.9999999999999998
* device instance $3 r0 *1 5.69,10.165 sg13_lv_pmos
M$3 \$6 \$4 \$1 \$6 sg13_lv_pmos W=1.1199999999999999 L=0.12999999999999995
* device instance $4 r0 *1 13.042,19.456 sg13_lv_pmos
M$4 vdda \$1 vout vdda sg13_lv_pmos W=0.9999999999999998 L=0.9999999999999998
* device instance $5 r0 *1 1.395,5.482 cap_cmim
C$5 \$1 vss cap_cmim w=7 l=7 m=1
.ENDS lvs_test

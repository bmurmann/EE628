* Extracted by KLayout with SG13G2 LVS runset on : 09/05/2024 10:00

* cell comp_5_split2
* pin sub!
.SUBCKT comp_5_split2 sub!
* device instance $1 r0 *1 -2.191,-4.403 sg13_lv_nmos
M$1 sub! \$2 \$3 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $2 r0 *1 -2.149,-0.904 sg13_lv_nmos
M$2 \$7 \$4 \$3 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $3 r0 *1 -3.449,-1.539 sg13_lv_pmos
M$3 \$7 \$2 \$8 \$8 sg13_lv_pmos W=4.0 L=0.13
* device instance $4 r0 *1 -0.007,-1.539 sg13_lv_pmos
M$4 \$8 \$4 \$7 \$8 sg13_lv_pmos W=4.0 L=0.13
.ENDS comp_5_split2

** sch_path: /foss/designs/Kate1/IDSM2.sch
**.subckt IDSM2 vhi vlo vdda vssa vin dout res clk
*.ipin vlo
*.ipin vdda
*.ipin vssa
*.ipin vin
*.ipin vhi
*.ipin res
*.ipin clk
*.opin dout
x1 res p1e p1 p2 vhi vdda vin vout1 vssa net3 net2 vlo stage_T6
x2 res p2e p2 p1 vhi vdda vout1 vout2 vssa vmid2 net1 vlo stage_T6
x4 p1e p1 clk p2 p2e clkgen_T6
x3 vdda p2 net1 vmid2 vssa net2 dout p1 vout2 res comparator_T6
**.ends

* expanding   symbol:  /foss/designs/Kate1/stage_T6.sym # of pins=12
** sym_path: /foss/designs/Kate1/stage_T6.sym
** sch_path: /foss/designs/Kate1/stage_T6.sch
.subckt stage_T6 res pse ps pr vhi vdda vin vout vssa vmid d vlo
*.iopin vhi
*.ipin pr
*.opin vout
*.ipin d
*.ipin vin
*.ipin ps
*.ipin pse
*.ipin res
*.opin vmid
*.iopin vlo
*.iopin vssa
*.iopin vdda
x1 pr d VDD VSS gn sg13g2_and2_1
x2 d pr VDD VSS gp sg13g2_nand2b_1
XC1 vx2 vx1 cap_cmim W=5.77e-6 L=5.77e-6 MF=1
XM3 vx1 psb vin vdda sg13_lv_pmos W=6.0u L=0.13u ng=3 m=1
XM4 vx1 ps vin vssa sg13_lv_nmos W=2.0u L=0.13u ng=1 m=1
XM5 vx1 gn vlo vssa sg13_lv_nmos W=0.5u L=0.13u ng=1 m=1
XM6 vx1 gp vhi vdda sg13_lv_pmos W=1.5u L=0.13u ng=1 m=1
XM7 vx2 pse vmid vssa sg13_lv_nmos W=2u L=0.13u ng=1 m=1
XM8 vx4 pr vx2 vssa sg13_lv_nmos W=2u L=0.13u ng=1 m=1
XC2 vx3 vx2 cap_cmim W=8.16e-6 L=8.16e-6 MF=1
XM9 vx4 ps vx3 vssa sg13_lv_nmos W=2u L=0.13u ng=1 m=1
XC3 vx4 vout cap_cmim W=8.16e-6 L=8.16e-6 MF=1
XM10 vout res vx4 vssa sg13_lv_nmos W=2u L=0.13u ng=1 m=1
XM11 vout vx3 vdda vdda sg13_lv_pmos W=10u L=1.5u ng=4 m=1
XM12 vout vx3 vssa vssa sg13_lv_nmos W=2.5u L=1.5u ng=1 m=1
XM1 vmid vmid vdda vdda sg13_lv_pmos W=10u L=1.5u ng=4 m=1
XM2 vmid vmid vssa vssa sg13_lv_nmos W=2.5u L=1.5u ng=1 m=1
x3 ps VDD VSS psb sg13g2_inv_1
.ends


* expanding   symbol:  /foss/designs/Kate1/clkgen_T6.sym # of pins=5
** sym_path: /foss/designs/Kate1/clkgen_T6.sym
** sch_path: /foss/designs/Kate1/clkgen_T6.sch
.subckt clkgen_T6 p1e p1 clkin p2 p2e
*.ipin clkin
*.opin p1e
*.opin p1
*.opin p2
*.opin p2e
x23 clkin VDD VSS clkinb sg13g2_inv_2
x2 clkinb VDD VSS clkinbb sg13g2_inv_2
x3 b1 clkinb VDD VSS net7 sg13g2_nand2_2
x4 clkinbb b2 VDD VSS net1 sg13g2_nand2_2
x14 net2 VDD VSS net3 sg13g2_inv_4
x1 net1 VDD VSS net2 sg13g2_inv_4
x5 net3 VDD VSS net4 sg13g2_inv_4
x6 net4 VDD VSS a1 sg13g2_inv_4
x7 a1 VDD VSS p1e sg13g2_inv_4
x8 p1e VDD VSS b1 sg13g2_inv_4
x9 p2e VDD VSS b2 sg13g2_inv_4
x10 a2 VDD VSS p2e sg13g2_inv_4
x15 net10 VDD VSS a2 sg13g2_inv_4
x16 net9 VDD VSS net10 sg13g2_inv_4
x17 net8 VDD VSS net9 sg13g2_inv_4
x18 net7 VDD VSS net8 sg13g2_inv_4
x11 a1 b1 VDD VSS net5 sg13g2_nand2_2
x19 a2 b2 VDD VSS net11 sg13g2_nand2_2
x12 net5 VDD VSS net6 sg13g2_inv_4
x20 net11 VDD VSS net12 sg13g2_inv_4
x13 net6 VDD VSS p1 sg13g2_inv_8
x21 net12 VDD VSS p2 sg13g2_inv_8
.ends


* expanding   symbol:  /foss/designs/Kate1/comparator_T6.sym # of pins=10
** sym_path: /foss/designs/Kate1/comparator_T6.sym
** sch_path: /foss/designs/Kate1/comparator_T6.sch
.subckt comparator_T6 vdda pc d vinp vssa dd dout ps vinm res
*.ipin pc
*.opin d
*.iopin vdda
*.ipin vinp
*.iopin vssa
*.ipin ps
*.ipin vinm
*.ipin res
*.opin dd
*.opin dout
x1 ps VDD VSS net5 sg13g2_inv_1
x2 din VDD VSS d sg13g2_buf_2
XC1 vinm_samp vssa cap_cmim W=5.77e-6 L=5.77e-6 MF=1
XM1 out1m pc vdda vdda sg13_lv_pmos W=4.0u L=0.13u ng=1 m=1
XM2 out1p out1m net3 vssa sg13_lv_nmos W=2.0u L=0.13u ng=1 m=1
XM3 out1m out1p vdda vdda sg13_lv_pmos W=4.0u L=0.13u ng=1 m=1
XM4 out1p out1m vdda vdda sg13_lv_pmos W=4.0u L=0.13u ng=1 m=1
XM5 out1p pc vdda vdda sg13_lv_pmos W=4.0u L=0.13u ng=1 m=1
XM6 out1m out1p net1 vssa sg13_lv_nmos W=2.0u L=0.13u ng=1 m=1
XM7 net3 pc net4 vssa sg13_lv_nmos W=2.0u L=0.13u ng=1 m=1
XM8 net1 pc net2 vssa sg13_lv_nmos W=2.0u L=0.13u ng=1 m=1
XM9 net4 vinm_samp vssa vssa sg13_lv_nmos W=2.0u L=1u ng=1 m=1
XM10 net2 vinp vssa vssa sg13_lv_nmos W=2.0u L=1u ng=1 m=1
XM11 vinm_samp net5 vinm vdda sg13_lv_pmos W=6.0u L=0.13u ng=3 m=1
XM12 vinm_samp ps vinm vssa sg13_lv_nmos W=2.0u L=0.13u ng=1 m=1
XM13 net6 out1p VDD VDD sg13_lv_pmos W=4.0u L=0.13u ng=1 m=1
XM14 din net6 net8 VSS sg13_lv_nmos W=2.0u L=0.13u ng=1 m=1
XM15 net6 din VDD VDD sg13_lv_pmos W=4.0u L=0.13u ng=1 m=1
XM16 din net6 VDD VDD sg13_lv_pmos W=4.0u L=0.13u ng=1 m=1
XM17 din out1m VDD VDD sg13_lv_pmos W=4.0u L=0.13u ng=1 m=1
XM18 net6 din net7 VSS sg13_lv_nmos W=2.0u L=0.13u ng=1 m=1
XM19 net8 out1m VSS VSS sg13_lv_nmos W=2.0u L=0.13u ng=1 m=1
XM20 net7 out1p VSS VSS sg13_lv_nmos W=2.0u L=0.13u ng=1 m=1
x4 res VDD VSS resb sg13g2_inv_1
x5 ps din dd net9 resb VDD VSS sg13g2_dfrbp_2
x3 dd VDD VSS dout sg13g2_inv_2
.ends

.GLOBAL VDD
.GLOBAL VSS
.end

* Extracted by KLayout with SG13G2 LVS runset on : 05/05/2024 06:21

* cell clock_5_split4
.SUBCKT clock_5_split4
* device instance $1 r0 *1 -0.448,0.074 sg13_lv_nmos
M$1 \$2 nand_B2 sub! sub! sg13_lv_nmos W=1.44 L=0.13
* device instance $3 r0 *1 0.582,0.074 sg13_lv_nmos
M$3 \$2 nand_A2 \$8 sub! sg13_lv_nmos W=1.44 L=0.13
* device instance $5 r0 *1 4.316,0.099 sg13_lv_nmos
M$5 sub! \$8 \$9 sub! sg13_lv_nmos W=2.96 L=0.13
* device instance $9 r0 *1 9.531,0.099 sg13_lv_nmos
M$9 sub! \$9 \$10 sub! sg13_lv_nmos W=2.96 L=0.13
* device instance $13 r0 *1 14.467,0.099 sg13_lv_nmos
M$13 sub! \$10 inv_bottom sub! sg13_lv_nmos W=2.96 L=0.13
* device instance $17 r0 *1 -0.448,1.759 sg13_lv_pmos
M$17 \$16 nand_B2 \$8 \$16 sg13_lv_pmos W=2.24 L=0.13
* device instance $19 r0 *1 0.582,1.759 sg13_lv_pmos
M$19 \$16 nand_A2 \$8 \$16 sg13_lv_pmos W=2.24 L=0.13
* device instance $21 r0 *1 4.316,1.759 sg13_lv_pmos
M$21 \$16 \$8 \$9 \$16 sg13_lv_pmos W=4.48 L=0.13
* device instance $25 r0 *1 9.531,1.759 sg13_lv_pmos
M$25 \$16 \$9 \$10 \$16 sg13_lv_pmos W=4.48 L=0.13
* device instance $29 r0 *1 14.467,1.759 sg13_lv_pmos
M$29 \$16 \$10 inv_bottom \$16 sg13_lv_pmos W=4.48 L=0.13
.ENDS clock_5_split4

* Extracted by KLayout with SG13G2 LVS runset on : 03/05/2024 04:44

* cell sg13g2_DCNDiode
* pin sub!
.SUBCKT sg13g2_DCNDiode sub!
* device instance $1 r0 *1 16.53,2.88 dantenna
D$1 sub! \$5 dantenna A=35.0028 P=58.08 m=1
* device instance $2 r0 *1 16.53,7.38 dantenna
D$2 sub! \$9 dantenna A=35.0028 P=58.08 m=1
.ENDS sg13g2_DCNDiode

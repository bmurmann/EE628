* Extracted by KLayout with SG13G2 LVS runset on : 06/05/2024 23:05

* cell UHEE628_S2024
* pin RES
* pin CK4
* pin CK5
* pin CK6
* pin IOVDD
* pin AVDD
* pin VDD
* pin IN6
* pin OUT6
* pin IN5
* pin OUT5
* pin IN4
* pin OUT4
* pin VLO
* pin VHI
* pin IN3
* pin OUT3
* pin VLDO
* pin IN2
* pin OUT2
* pin IN1
* pin OUT1
* pin VREF
* pin CK3
* pin CK2
* pin CK1
* pin VSS
.SUBCKT UHEE628_S2024 RES CK4 CK5 CK6 IOVDD AVDD VDD IN6 OUT6 IN5 OUT5 IN4 OUT4
+ VLO VHI IN3 OUT3 VLDO IN2 OUT2 IN1 OUT1 VREF CK3 CK2 CK1 VSS
* device instance $1 r0 *1 500.255,239.005 sg13_lv_nmos
M$1 \$181 \$186 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $2 r0 *1 700.255,239.005 sg13_lv_nmos
M$2 \$182 \$187 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $3 r0 *1 800.255,239.005 sg13_lv_nmos
M$3 \$183 \$188 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $4 r0 *1 900.255,239.005 sg13_lv_nmos
M$4 \$184 \$189 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $5 r0 *1 1060.995,297.48 sg13_lv_nmos
M$5 \$235 \$237 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $6 r0 *1 1060.995,300.99 sg13_lv_nmos
M$6 \$263 \$237 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $7 r0 *1 1060.995,397.48 sg13_lv_nmos
M$7 \$350 \$352 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $8 r0 *1 1060.995,400.99 sg13_lv_nmos
M$8 \$378 \$352 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $9 r0 *1 1060.995,497.48 sg13_lv_nmos
M$9 \$465 \$467 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $10 r0 *1 1060.995,500.99 sg13_lv_nmos
M$10 \$493 \$467 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $11 r0 *1 485.618,504.427 sg13_lv_nmos
M$11 \$517 \$527 \$533 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $12 r0 *1 486.008,504.427 sg13_lv_nmos
M$12 \$533 \$518 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $13 r0 *1 486.568,504.427 sg13_lv_nmos
M$13 VSS \$504 \$532 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $14 r0 *1 486.923,504.427 sg13_lv_nmos
M$14 \$532 \$517 \$518 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $15 r0 *1 483.978,504.537 sg13_lv_nmos
M$15 VSS \$515 \$516 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $16 r0 *1 484.648,504.537 sg13_lv_nmos
M$16 \$516 \$510 \$517 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $17 r0 *1 482.098,504.652 sg13_lv_nmos
M$17 \$514 \$527 \$515 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $18 r0 *1 482.608,504.652 sg13_lv_nmos
M$18 \$515 \$510 \$531 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $19 r0 *1 482.998,504.652 sg13_lv_nmos
M$19 \$531 \$516 \$530 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $20 r0 *1 483.358,504.652 sg13_lv_nmos
M$20 VSS \$504 \$530 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $21 r0 *1 476.768,504.592 sg13_lv_nmos
M$21 VSS \$689 \$513 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $22 r0 *1 487.963,504.592 sg13_lv_nmos
M$22 VSS \$517 \$519 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $23 r0 *1 489.163,504.497 sg13_lv_nmos
M$23 \$520 \$517 VSS VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $24 r0 *1 489.703,504.592 sg13_lv_nmos
M$24 VSS \$520 \$521 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $25 r0 *1 491.898,504.592 sg13_lv_nmos
M$25 VSS \$521 \$467 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $27 r0 *1 494.693,504.591 sg13_lv_nmos
M$27 VSS \$181 \$504 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $28 r0 *1 496.608,504.591 sg13_lv_nmos
M$28 VSS \$534 \$522 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $30 r0 *1 497.628,504.641 sg13_lv_nmos
M$30 VSS \$584 \$534 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $31 r0 *1 478.818,504.452 sg13_lv_nmos
M$31 \$514 \$584 \$529 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $32 r0 *1 479.188,504.452 sg13_lv_nmos
M$32 \$529 \$504 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $33 r0 *1 480.333,504.767 sg13_lv_nmos
M$33 VSS \$689 \$527 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $34 r0 *1 480.843,504.767 sg13_lv_nmos
M$34 VSS \$527 \$510 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $35 r0 *1 481.503,510.997 sg13_lv_nmos
M$35 VSS \$569 \$574 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $36 r0 *1 481.703,513.099 sg13_lv_nmos
M$36 \$574 \$631 \$580 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $37 r0 *1 483.503,509.467 sg13_lv_nmos
M$37 \$564 \$689 \$565 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $38 r0 *1 482.903,513.099 sg13_lv_nmos
M$38 \$580 \$600 \$581 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $39 r0 *1 484.103,513.099 sg13_lv_nmos
M$39 \$600 \$581 \$582 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $40 r0 *1 485.503,510.997 sg13_lv_nmos
M$40 VSS \$565 \$575 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $41 r0 *1 485.303,513.099 sg13_lv_nmos
M$41 \$582 \$631 \$575 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $42 r0 *1 488.561,513.099 sg13_lv_nmos
M$42 VSS \$600 \$583 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $43 r0 *1 489.761,513.099 sg13_lv_nmos
M$43 \$583 \$584 \$609 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $44 r0 *1 490.961,513.099 sg13_lv_nmos
M$44 \$584 \$609 \$585 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $45 r0 *1 492.161,513.099 sg13_lv_nmos
M$45 \$585 \$581 VSS VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $46 r0 *1 438.155,518.846 sg13_lv_nmos
M$46 VSS \$622 \$623 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $50 r0 *1 441.035,518.846 sg13_lv_nmos
M$50 VSS \$623 \$624 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $54 r0 *1 443.915,518.846 sg13_lv_nmos
M$54 VSS \$624 \$625 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $58 r0 *1 446.795,518.846 sg13_lv_nmos
M$58 VSS \$625 \$626 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $62 r0 *1 449.675,518.846 sg13_lv_nmos
M$62 VSS \$626 \$627 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $66 r0 *1 452.555,518.846 sg13_lv_nmos
M$66 VSS \$627 \$628 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $70 r0 *1 458.315,518.846 sg13_lv_nmos
M$70 VSS \$629 \$630 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $74 r0 *1 461.135,518.846 sg13_lv_nmos
M$74 VSS \$630 \$631 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $82 r0 *1 431.455,521.281 sg13_lv_nmos
M$82 VSS \$182 \$633 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $84 r0 *1 433.375,521.281 sg13_lv_nmos
M$84 VSS \$633 \$679 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $86 r0 *1 435.35,518.871 sg13_lv_nmos
M$86 \$657 \$686 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $88 r0 *1 436.38,518.871 sg13_lv_nmos
M$88 \$657 \$633 \$622 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $90 r0 *1 435.35,521.256 sg13_lv_nmos
M$90 \$680 \$628 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $92 r0 *1 436.38,521.256 sg13_lv_nmos
M$92 \$680 \$679 \$707 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $94 r0 *1 438.155,521.281 sg13_lv_nmos
M$94 VSS \$707 \$681 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $98 r0 *1 441.035,521.281 sg13_lv_nmos
M$98 VSS \$681 \$682 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $102 r0 *1 443.915,521.281 sg13_lv_nmos
M$102 VSS \$682 \$683 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $106 r0 *1 446.795,521.281 sg13_lv_nmos
M$106 VSS \$683 \$684 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $110 r0 *1 449.675,521.281 sg13_lv_nmos
M$110 VSS \$684 \$685 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $114 r0 *1 452.555,521.281 sg13_lv_nmos
M$114 VSS \$685 \$686 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $118 r0 *1 455.51,518.871 sg13_lv_nmos
M$118 \$658 \$628 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $120 r0 *1 456.54,518.871 sg13_lv_nmos
M$120 \$658 \$626 \$629 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $122 r0 *1 455.51,521.256 sg13_lv_nmos
M$122 \$687 \$686 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $124 r0 *1 456.54,521.256 sg13_lv_nmos
M$124 \$687 \$684 \$692 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $126 r0 *1 458.315,521.281 sg13_lv_nmos
M$126 VSS \$692 \$688 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $130 r0 *1 461.135,521.281 sg13_lv_nmos
M$130 VSS \$688 \$689 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $138 r0 *1 431.5,535.261 sg13_lv_nmos
M$138 VSS \$689 \$731 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $139 r0 *1 432.935,535.356 sg13_lv_nmos
M$139 VSS \$521 \$732 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $140 r0 *1 433.785,535.261 sg13_lv_nmos
M$140 VSS \$631 \$750 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $141 r0 *1 434.095,535.261 sg13_lv_nmos
M$141 \$750 \$732 \$733 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $142 r0 *1 434.07,553.206 sg13_lv_nmos
M$142 \$791 \$735 VLO VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $143 r0 *1 435.785,535.421 sg13_lv_nmos
M$143 \$734 \$631 \$747 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $144 r0 *1 436.295,535.421 sg13_lv_nmos
M$144 VSS \$521 \$747 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $145 r0 *1 436.805,535.371 sg13_lv_nmos
M$145 VSS \$734 \$735 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $146 r0 *1 436.815,553.216 sg13_lv_nmos
M$146 \$791 \$689 \$587 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $147 r0 *1 443.55,535.276 sg13_lv_nmos
M$147 VSS \$736 \$736 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $148 r0 *1 444.09,553.171 sg13_lv_nmos
M$148 \$736 \$685 \$789 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $149 r0 *1 449.83,597.155 sg13_lv_nmos
M$149 \$857 \$910 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $151 r0 *1 450.86,597.155 sg13_lv_nmos
M$151 \$857 \$867 \$868 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $153 r0 *1 455.2,535.261 sg13_lv_nmos
M$153 VSS \$757 \$752 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $154 r0 *1 454.14,553.166 sg13_lv_nmos
M$154 \$789 \$631 \$797 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $155 r0 *1 455.45,553.166 sg13_lv_nmos
M$155 \$797 \$689 \$757 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $156 r0 *1 456.763,553.166 sg13_lv_nmos
M$156 \$797 \$181 \$752 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $157 r0 *1 466.5,535.261 sg13_lv_nmos
M$157 VSS \$631 \$737 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $158 r0 *1 467.935,535.356 sg13_lv_nmos
M$158 VSS \$522 \$738 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $159 r0 *1 468.785,535.261 sg13_lv_nmos
M$159 VSS \$689 \$745 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $160 r0 *1 469.095,535.261 sg13_lv_nmos
M$160 \$745 \$738 \$739 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $161 r0 *1 469.07,553.206 sg13_lv_nmos
M$161 \$792 \$741 VLO VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $162 r0 *1 469.99,597.155 sg13_lv_nmos
M$162 \$864 \$863 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $164 r0 *1 471.02,597.155 sg13_lv_nmos
M$164 \$864 \$861 \$869 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $166 r0 *1 470.785,535.421 sg13_lv_nmos
M$166 \$740 \$689 \$743 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $167 r0 *1 471.295,535.421 sg13_lv_nmos
M$167 VSS \$522 \$743 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $168 r0 *1 471.805,535.371 sg13_lv_nmos
M$168 VSS \$740 \$741 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $169 r0 *1 471.815,553.216 sg13_lv_nmos
M$169 \$792 \$631 \$752 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $170 r0 *1 478.55,535.276 sg13_lv_nmos
M$170 VSS \$569 \$569 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $171 r0 *1 479.09,553.171 sg13_lv_nmos
M$171 \$569 \$627 \$790 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $172 r0 *1 490.2,535.261 sg13_lv_nmos
M$172 VSS \$758 \$564 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $173 r0 *1 489.14,553.166 sg13_lv_nmos
M$173 \$790 \$689 \$798 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $174 r0 *1 490.45,553.166 sg13_lv_nmos
M$174 \$798 \$631 \$758 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $175 r0 *1 491.763,553.166 sg13_lv_nmos
M$175 \$798 \$181 \$564 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $176 r0 *1 452.635,597.18 sg13_lv_nmos
M$176 VSS \$868 \$858 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $180 r0 *1 455.515,597.18 sg13_lv_nmos
M$180 VSS \$858 \$859 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $184 r0 *1 458.395,597.18 sg13_lv_nmos
M$184 VSS \$859 \$860 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $188 r0 *1 461.275,597.18 sg13_lv_nmos
M$188 VSS \$860 \$861 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $192 r0 *1 464.155,597.18 sg13_lv_nmos
M$192 VSS \$861 \$862 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $196 r0 *1 467.035,597.18 sg13_lv_nmos
M$196 VSS \$862 \$863 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $200 r0 *1 472.795,597.18 sg13_lv_nmos
M$200 VSS \$869 \$865 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $204 r0 *1 475.615,597.18 sg13_lv_nmos
M$204 VSS \$865 \$866 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $212 r0 *1 445.935,602.98 sg13_lv_nmos
M$212 VSS \$853 \$867 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $214 r0 *1 447.855,602.98 sg13_lv_nmos
M$214 VSS \$867 \$903 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $216 r0 *1 449.83,602.955 sg13_lv_nmos
M$216 \$904 \$863 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $218 r0 *1 450.86,602.955 sg13_lv_nmos
M$218 \$904 \$903 \$914 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $220 r0 *1 452.635,602.98 sg13_lv_nmos
M$220 VSS \$914 \$905 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $224 r0 *1 455.515,602.98 sg13_lv_nmos
M$224 VSS \$905 \$906 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $228 r0 *1 458.395,602.98 sg13_lv_nmos
M$228 VSS \$906 \$907 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $232 r0 *1 461.275,602.98 sg13_lv_nmos
M$232 VSS \$907 \$908 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $236 r0 *1 464.155,602.98 sg13_lv_nmos
M$236 VSS \$908 \$909 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $240 r0 *1 467.035,602.98 sg13_lv_nmos
M$240 VSS \$909 \$910 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $244 r0 *1 469.99,602.955 sg13_lv_nmos
M$244 \$911 \$910 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $246 r0 *1 471.02,602.955 sg13_lv_nmos
M$246 \$911 \$908 \$915 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $248 r0 *1 472.795,602.98 sg13_lv_nmos
M$248 VSS \$915 \$912 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $252 r0 *1 475.615,602.98 sg13_lv_nmos
M$252 VSS \$912 \$913 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $260 r0 *1 433.27,616.415 sg13_lv_nmos
M$260 VSS \$913 \$975 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $261 r0 *1 434.36,616.51 sg13_lv_nmos
M$261 VSS \$946 \$979 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $262 r0 *1 435.21,616.415 sg13_lv_nmos
M$262 VSS \$866 \$988 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $263 r0 *1 435.52,616.415 sg13_lv_nmos
M$263 \$988 \$979 \$976 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $264 r0 *1 436.85,616.575 sg13_lv_nmos
M$264 \$984 \$866 \$996 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $265 r0 *1 437.36,616.575 sg13_lv_nmos
M$265 VSS \$946 \$996 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $266 r0 *1 437.87,616.525 sg13_lv_nmos
M$266 VSS \$984 \$967 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $267 r0 *1 441.655,618.475 sg13_lv_nmos
M$267 VLO \$967 \$1015 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $268 r0 *1 454.37,616.04 sg13_lv_nmos
M$268 \$968 \$909 \$993 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $269 r0 *1 454.37,616.55 sg13_lv_nmos
M$269 \$993 \$866 \$1071 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $270 r0 *1 454.37,617.83 sg13_lv_nmos
M$270 \$1105 \$913 \$1071 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $271 r0 *1 454.37,618.34 sg13_lv_nmos
M$271 \$1071 \$181 \$1016 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $272 r0 *1 469.325,616.415 sg13_lv_nmos
M$272 VSS \$866 \$977 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $273 r0 *1 470.415,616.51 sg13_lv_nmos
M$273 VSS \$947 \$980 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $274 r0 *1 471.265,616.415 sg13_lv_nmos
M$274 VSS \$913 \$991 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $275 r0 *1 471.575,616.415 sg13_lv_nmos
M$275 \$991 \$980 \$978 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $276 r0 *1 472.905,616.575 sg13_lv_nmos
M$276 \$985 \$913 \$1004 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $277 r0 *1 473.415,616.575 sg13_lv_nmos
M$277 VSS \$947 \$1004 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $278 r0 *1 473.925,616.525 sg13_lv_nmos
M$278 VSS \$985 \$969 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $279 r0 *1 477.71,618.475 sg13_lv_nmos
M$279 VLO \$969 \$1017 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $280 r0 *1 490.425,617.83 sg13_lv_nmos
M$280 \$1106 \$866 \$1072 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $281 r0 *1 490.425,618.34 sg13_lv_nmos
M$281 \$1072 \$181 \$1018 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $282 r0 *1 490.425,616.04 sg13_lv_nmos
M$282 \$970 \$862 \$994 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $283 r0 *1 490.425,616.55 sg13_lv_nmos
M$283 \$994 \$913 \$1072 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $284 r0 *1 505.425,616.53 sg13_lv_nmos
M$284 VSS \$913 \$981 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $285 r0 *1 520.915,619.83 sg13_lv_nmos
M$285 \$1037 \$1047 \$1049 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $286 r0 *1 521.225,619.83 sg13_lv_nmos
M$286 \$1049 \$1033 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $287 r0 *1 521.805,620.215 sg13_lv_nmos
M$287 VSS \$1062 \$1038 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $288 r0 *1 522.895,619.895 sg13_lv_nmos
M$288 VSS \$1033 \$1050 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $289 r0 *1 523.205,619.895 sg13_lv_nmos
M$289 \$1050 \$1038 \$1046 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $290 r0 *1 528.06,620.215 sg13_lv_nmos
M$290 \$1048 \$1039 \$1040 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $291 r0 *1 528.595,620.055 sg13_lv_nmos
M$291 \$1038 \$1073 \$1048 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $292 r0 *1 529.645,619.83 sg13_lv_nmos
M$292 \$1040 \$1041 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $293 r0 *1 530.155,619.83 sg13_lv_nmos
M$293 VSS \$1033 \$1052 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $294 r0 *1 530.465,619.83 sg13_lv_nmos
M$294 \$1052 \$1048 \$1041 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $295 r0 *1 532.505,619.94 sg13_lv_nmos
M$295 VSS \$1048 \$1043 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $296 r0 *1 531.485,619.99 sg13_lv_nmos
M$296 VSS \$1048 \$1042 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $298 r0 *1 533.525,619.99 sg13_lv_nmos
M$298 VSS \$1043 \$946 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $300 r0 *1 535.21,620.01 sg13_lv_nmos
M$300 VSS \$946 \$1010 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $302 r0 *1 537,620.005 sg13_lv_nmos
M$302 \$1033 \$181 VSS VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $303 r0 *1 433.495,621.675 sg13_lv_nmos
M$303 \$1344 \$913 \$1015 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $304 r0 *1 456.64,623.065 sg13_lv_nmos
M$304 VSS \$1105 \$1016 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $305 r0 *1 462.64,623.065 sg13_lv_nmos
M$305 VSS \$968 \$968 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $306 r0 *1 469.55,621.675 sg13_lv_nmos
M$306 \$1016 \$866 \$1017 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $307 r0 *1 492.695,623.065 sg13_lv_nmos
M$307 VSS \$1106 \$1018 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $308 r0 *1 498.695,623.065 sg13_lv_nmos
M$308 VSS \$970 \$970 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $309 r0 *1 505.05,623.5 sg13_lv_nmos
M$309 \$1061 \$913 \$1018 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $310 r0 *1 509.96,626.51 sg13_lv_nmos
M$310 VSS \$970 \$1115 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $311 r0 *1 514.885,626.51 sg13_lv_nmos
M$311 VSS \$1061 \$1116 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $312 r0 *1 523.98,620.62 sg13_lv_nmos
M$312 \$1037 \$1039 \$1062 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $313 r0 *1 524.49,620.62 sg13_lv_nmos
M$313 \$1062 \$1073 \$1046 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $314 r0 *1 525.75,620.095 sg13_lv_nmos
M$314 VSS \$1039 \$1073 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $315 r0 *1 526.85,620.095 sg13_lv_nmos
M$315 VSS \$913 \$1039 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $316 r0 *1 532.795,625.47 sg13_lv_nmos
M$316 VSS \$1103 \$947 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $318 r0 *1 532.845,626.49 sg13_lv_nmos
M$318 VSS \$1047 \$1103 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $319 r0 *1 522.75,627.29 sg13_lv_nmos
M$319 VSS \$1134 \$1117 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $320 r0 *1 529.69,627.28 sg13_lv_nmos
M$320 VSS \$1133 \$1118 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $321 r0 *1 509.855,627.99 sg13_lv_nmos
M$321 \$1115 \$866 \$1123 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $322 r0 *1 514.795,627.99 sg13_lv_nmos
M$322 \$1116 \$866 \$1124 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $323 r0 *1 523.03,628.795 sg13_lv_nmos
M$323 \$1117 \$1047 \$1129 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $324 r0 *1 529.34,628.76 sg13_lv_nmos
M$324 \$1118 \$1129 \$1047 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $325 r0 *1 509.835,629.77 sg13_lv_nmos
M$325 \$1123 \$1134 \$1133 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $326 r0 *1 514.62,629.77 sg13_lv_nmos
M$326 \$1124 \$1133 \$1134 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $327 r0 *1 1060.995,797.48 sg13_lv_nmos
M$327 \$1292 \$1010 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $328 r0 *1 1060.995,800.99 sg13_lv_nmos
M$328 \$1319 \$1010 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $329 r0 *1 633.21,835.705 sg13_lv_nmos
M$329 VSS \$1380 \$1380 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $331 r0 *1 630.06,842.755 sg13_lv_nmos
M$331 \$1391 \$1434 \$1384 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $333 r0 *1 622.76,843.455 sg13_lv_nmos
M$333 VSS \$1380 \$1396 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $335 r0 *1 626.34,843.455 sg13_lv_nmos
M$335 VSS \$1384 \$1397 VSS sg13_lv_nmos W=2.0 L=1.0
* device instance $337 r0 *1 623.505,845.055 sg13_lv_nmos
M$337 \$1396 \$1457 \$1402 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $339 r0 *1 626.465,845.055 sg13_lv_nmos
M$339 \$1397 \$1457 \$1403 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $341 r0 *1 632.73,845.055 sg13_lv_nmos
M$341 VSS \$1412 \$1404 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $343 r0 *1 635.69,845.055 sg13_lv_nmos
M$343 VSS \$1413 \$1405 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $345 r0 *1 592.87,846.075 sg13_lv_nmos
M$345 VSS \$1386 \$1406 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $347 r0 *1 614.46,846.075 sg13_lv_nmos
M$347 VSS \$1387 \$1391 VSS sg13_lv_nmos W=2.5 L=1.5
* device instance $349 r0 *1 623.505,846.655 sg13_lv_nmos
M$349 \$1402 \$1412 \$1413 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $351 r0 *1 626.465,846.655 sg13_lv_nmos
M$351 \$1403 \$1413 \$1412 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $353 r0 *1 632.73,846.655 sg13_lv_nmos
M$353 \$1404 \$1414 \$1419 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $355 r0 *1 635.69,846.655 sg13_lv_nmos
M$355 \$1405 \$1419 \$1414 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $357 r0 *1 585.345,846.95 sg13_lv_nmos
M$357 \$1417 \$1434 \$1854 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $359 r0 *1 586.14,851.955 sg13_lv_nmos
M$359 VLO \$1504 \$1417 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $360 r0 *1 588.475,849.383 sg13_lv_nmos
M$360 \$1382 \$1457 \$1420 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $361 r0 *1 588.475,852.473 sg13_lv_nmos
M$361 \$1382 \$1434 \$1386 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $362 r0 *1 589.55,849.383 sg13_lv_nmos
M$362 \$1420 \$1675 \$1380 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $363 r0 *1 606.935,846.95 sg13_lv_nmos
M$363 \$1418 \$1457 \$1406 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $365 r0 *1 607.73,851.955 sg13_lv_nmos
M$365 VLO \$1505 \$1418 VSS sg13_lv_nmos W=0.5 L=0.13
* device instance $366 r0 *1 610.065,849.383 sg13_lv_nmos
M$366 \$1383 \$1434 \$1421 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $367 r0 *1 610.065,852.473 sg13_lv_nmos
M$367 \$1383 \$1457 \$1387 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $368 r0 *1 611.14,849.383 sg13_lv_nmos
M$368 \$1421 \$1458 \$1380 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $369 r0 *1 623.635,852.165 sg13_lv_nmos
M$369 \$1490 \$1414 \$1523 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $370 r0 *1 623.945,852.165 sg13_lv_nmos
M$370 \$1523 \$1489 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $371 r0 *1 624.525,852.55 sg13_lv_nmos
M$371 VSS \$1535 \$1491 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $372 r0 *1 632.365,852.165 sg13_lv_nmos
M$372 \$1494 \$1495 VSS VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $373 r0 *1 632.875,852.165 sg13_lv_nmos
M$373 VSS \$1489 \$1528 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $374 r0 *1 633.185,852.165 sg13_lv_nmos
M$374 \$1528 \$1507 \$1495 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $375 r0 *1 635.225,852.275 sg13_lv_nmos
M$375 VSS \$1507 \$1497 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $376 r0 *1 634.205,852.325 sg13_lv_nmos
M$376 VSS \$1507 \$1496 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $378 r0 *1 636.245,852.325 sg13_lv_nmos
M$378 VSS \$1497 \$1590 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $380 r0 *1 620.94,852.345 sg13_lv_nmos
M$380 VSS \$1434 \$1422 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $381 r0 *1 622.38,852.345 sg13_lv_nmos
M$381 VSS \$181 \$1489 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $382 r0 *1 625.615,852.23 sg13_lv_nmos
M$382 VSS \$1489 \$1524 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $383 r0 *1 625.925,852.23 sg13_lv_nmos
M$383 \$1524 \$1491 \$1492 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $384 r0 *1 626.7,852.955 sg13_lv_nmos
M$384 \$1490 \$1493 \$1535 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $385 r0 *1 627.21,852.955 sg13_lv_nmos
M$385 \$1535 \$1506 \$1492 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $386 r0 *1 628.47,852.43 sg13_lv_nmos
M$386 VSS \$1493 \$1506 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $387 r0 *1 629.57,852.43 sg13_lv_nmos
M$387 VSS \$1434 \$1493 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $388 r0 *1 630.78,852.55 sg13_lv_nmos
M$388 \$1507 \$1493 \$1494 VSS sg13_lv_nmos W=0.42 L=0.13
* device instance $389 r0 *1 631.315,852.39 sg13_lv_nmos
M$389 \$1491 \$1506 \$1507 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $390 r0 *1 637.86,852.395 sg13_lv_nmos
M$390 VSS \$1414 \$1498 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $391 r0 *1 638.37,852.345 sg13_lv_nmos
M$391 VSS \$1498 \$1591 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $393 r0 *1 640.4,852.345 sg13_lv_nmos
M$393 VSS \$1590 \$1499 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $395 r0 *1 594.145,854.805 sg13_lv_nmos
M$395 \$1382 \$181 \$1406 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $399 r0 *1 615.735,854.805 sg13_lv_nmos
M$399 \$1383 \$181 \$1391 VSS sg13_lv_nmos W=2.0 L=0.13
* device instance $403 r0 *1 617.465,863.425 sg13_lv_nmos
M$403 \$1592 \$1626 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $405 r0 *1 618.495,863.425 sg13_lv_nmos
M$405 \$1592 \$1627 \$1607 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $407 r0 *1 640.7,863.425 sg13_lv_nmos
M$407 \$1598 \$1597 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $409 r0 *1 641.73,863.425 sg13_lv_nmos
M$409 \$1598 \$1596 \$1608 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $411 r0 *1 623.374,863.452 sg13_lv_nmos
M$411 VSS \$1593 \$1594 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $415 r0 *1 626.254,863.452 sg13_lv_nmos
M$415 VSS \$1594 \$1595 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $419 r0 *1 629.134,863.452 sg13_lv_nmos
M$419 VSS \$1595 \$1596 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $423 r0 *1 632.714,863.452 sg13_lv_nmos
M$423 VSS \$1596 \$1458 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $427 r0 *1 636.294,863.452 sg13_lv_nmos
M$427 VSS \$1458 \$1597 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $431 r0 *1 643.75,863.45 sg13_lv_nmos
M$431 VSS \$1608 \$1599 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $435 r0 *1 646.57,863.452 sg13_lv_nmos
M$435 VSS \$1599 \$1457 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $443 r0 *1 577.495,864.355 sg13_lv_nmos
M$443 \$1622 \$1457 \$1637 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $444 r0 *1 578.005,864.355 sg13_lv_nmos
M$444 VSS \$1590 \$1637 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $445 r0 *1 578.515,864.305 sg13_lv_nmos
M$445 VSS \$1622 \$1504 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $446 r0 *1 579.805,864.29 sg13_lv_nmos
M$446 VSS \$1590 \$1623 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $447 r0 *1 580.655,864.195 sg13_lv_nmos
M$447 VSS \$1457 \$1635 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $448 r0 *1 580.965,864.195 sg13_lv_nmos
M$448 \$1635 \$1623 \$1533 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $449 r0 *1 582.555,864.195 sg13_lv_nmos
M$449 VSS \$1434 \$1473 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $450 r0 *1 599.085,864.355 sg13_lv_nmos
M$450 \$1624 \$1434 \$1632 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $451 r0 *1 599.595,864.355 sg13_lv_nmos
M$451 VSS \$1591 \$1632 VSS sg13_lv_nmos W=0.64 L=0.13
* device instance $452 r0 *1 600.105,864.305 sg13_lv_nmos
M$452 VSS \$1624 \$1505 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $453 r0 *1 601.395,864.29 sg13_lv_nmos
M$453 VSS \$1591 \$1625 VSS sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $454 r0 *1 602.245,864.195 sg13_lv_nmos
M$454 VSS \$1434 \$1629 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $455 r0 *1 602.555,864.195 sg13_lv_nmos
M$455 \$1629 \$1625 \$1534 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $456 r0 *1 604.145,864.195 sg13_lv_nmos
M$456 VSS \$1457 \$1474 VSS sg13_lv_nmos W=0.74 L=0.13
* device instance $457 r0 *1 617.465,869.102 sg13_lv_nmos
M$457 \$1670 \$1597 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $459 r0 *1 618.495,869.102 sg13_lv_nmos
M$459 \$1670 \$1669 \$1678 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $461 r0 *1 620.494,869.122 sg13_lv_nmos
M$461 VSS \$1678 \$1671 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $465 r0 *1 620.494,863.454 sg13_lv_nmos
M$465 VSS \$1607 \$1593 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $469 r0 *1 623.374,869.122 sg13_lv_nmos
M$469 VSS \$1671 \$1672 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $473 r0 *1 626.254,869.122 sg13_lv_nmos
M$473 VSS \$1672 \$1673 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $477 r0 *1 629.134,869.122 sg13_lv_nmos
M$477 VSS \$1673 \$1674 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $481 r0 *1 632.714,869.122 sg13_lv_nmos
M$481 VSS \$1674 \$1675 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $485 r0 *1 636.294,869.122 sg13_lv_nmos
M$485 VSS \$1675 \$1626 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $489 r0 *1 640.44,869.102 sg13_lv_nmos
M$489 \$1676 \$1626 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $491 r0 *1 641.47,869.102 sg13_lv_nmos
M$491 \$1676 \$1674 \$1679 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $493 r0 *1 643.505,869.122 sg13_lv_nmos
M$493 VSS \$1679 \$1677 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $497 r0 *1 613.57,869.127 sg13_lv_nmos
M$497 VSS \$1692 \$1627 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $499 r0 *1 615.49,869.127 sg13_lv_nmos
M$499 VSS \$1627 \$1669 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $501 r0 *1 646.325,869.128 sg13_lv_nmos
M$501 VSS \$1677 \$1434 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $509 r0 *1 1060.995,897.48 sg13_lv_nmos
M$509 \$1802 \$1499 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $510 r0 *1 1060.995,900.99 sg13_lv_nmos
M$510 \$1829 \$1499 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $511 r0 *1 1060.995,997.48 sg13_lv_nmos
M$511 \$1916 \$1924 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $512 r0 *1 1060.995,1000.99 sg13_lv_nmos
M$512 \$1944 \$1924 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $513 r0 *1 700.255,1060.995 sg13_lv_nmos
M$513 \$853 \$2010 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $514 r0 *1 800.255,1060.995 sg13_lv_nmos
M$514 \$1692 \$2011 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $515 r0 *1 900.255,1060.995 sg13_lv_nmos
M$515 \$2005 \$2012 VSS VSS sg13_lv_nmos W=2.75 L=0.13
* device instance $516 r0 *1 501.765,239.055 sg13_hv_nmos
M$516 VSS \$129 \$186 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $517 r0 *1 701.765,239.055 sg13_hv_nmos
M$517 VSS \$130 \$187 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $518 r0 *1 801.765,239.055 sg13_hv_nmos
M$518 VSS \$132 \$188 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $519 r0 *1 901.765,239.055 sg13_hv_nmos
M$519 VSS \$133 \$189 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $520 r0 *1 90.95,285.52 sg13_hv_nmos
M$520 VSS \$225 IN6 VSS sg13_hv_nmos W=88.00000000000001 L=0.5999999999999999
* device instance $540 r0 *1 1209.05,294.58 sg13_hv_nmos
M$540 VSS \$252 OUT6 VSS sg13_hv_nmos W=35.199999999999996 L=0.5999999999999999
* device instance $548 r0 *1 1064.68,297.64 sg13_hv_nmos
M$548 \$236 \$237 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $549 r0 *1 1064.68,298.47 sg13_hv_nmos
M$549 VSS \$235 \$246 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $550 r0 *1 1064.68,299.81 sg13_hv_nmos
M$550 VSS \$246 \$252 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $551 r0 *1 1064.68,301.15 sg13_hv_nmos
M$551 \$264 \$237 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $552 r0 *1 1064.68,301.98 sg13_hv_nmos
M$552 VSS \$263 \$271 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $553 r0 *1 1064.68,303.32 sg13_hv_nmos
M$553 VSS \$271 \$216 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $554 r0 *1 90.95,385.52 sg13_hv_nmos
M$554 VSS \$340 IN5 VSS sg13_hv_nmos W=88.00000000000001 L=0.5999999999999999
* device instance $574 r0 *1 1209.05,394.58 sg13_hv_nmos
M$574 VSS \$367 OUT5 VSS sg13_hv_nmos W=35.199999999999996 L=0.5999999999999999
* device instance $582 r0 *1 1064.68,397.64 sg13_hv_nmos
M$582 \$351 \$352 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $583 r0 *1 1064.68,398.47 sg13_hv_nmos
M$583 VSS \$350 \$361 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $584 r0 *1 1064.68,399.81 sg13_hv_nmos
M$584 VSS \$361 \$367 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $585 r0 *1 1064.68,401.15 sg13_hv_nmos
M$585 \$379 \$352 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $586 r0 *1 1064.68,401.98 sg13_hv_nmos
M$586 VSS \$378 \$386 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $587 r0 *1 1064.68,403.32 sg13_hv_nmos
M$587 VSS \$386 \$331 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $588 r0 *1 90.95,485.52 sg13_hv_nmos
M$588 VSS \$455 IN4 VSS sg13_hv_nmos W=88.00000000000001 L=0.5999999999999999
* device instance $608 r0 *1 1209.05,494.58 sg13_hv_nmos
M$608 VSS \$482 OUT4 VSS sg13_hv_nmos W=35.199999999999996 L=0.5999999999999999
* device instance $616 r0 *1 1064.68,497.64 sg13_hv_nmos
M$616 \$466 \$467 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $617 r0 *1 1064.68,498.47 sg13_hv_nmos
M$617 VSS \$465 \$476 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $618 r0 *1 1064.68,499.81 sg13_hv_nmos
M$618 VSS \$476 \$482 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $619 r0 *1 1064.68,501.15 sg13_hv_nmos
M$619 \$494 \$467 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $620 r0 *1 1064.68,501.98 sg13_hv_nmos
M$620 VSS \$493 \$501 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $621 r0 *1 1064.68,503.32 sg13_hv_nmos
M$621 VSS \$501 \$446 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $622 r0 *1 90.95,585.52 sg13_hv_nmos
M$622 VSS \$845 VLO VSS sg13_hv_nmos W=88.00000000000001 L=0.5999999999999999
* device instance $642 r0 *1 1139.21,663.22 sg13_hv_nmos
M$642 VSS \$1185 \$1184 VSS sg13_hv_nmos W=108.0 L=0.5
* device instance $648 r0 *1 1139.21,673 sg13_hv_nmos
M$648 VSS \$1185 VSS VSS sg13_hv_nmos W=126.0 L=9.5
* device instance $668 r0 *1 1194.53,668.155 sg13_hv_nmos
M$668 VSS \$1184 IOVDD VSS sg13_hv_nmos W=756.7999999999977 L=0.5999999999999999
* device instance $840 r0 *1 90.95,685.52 sg13_hv_nmos
M$840 VSS \$1190 VHI VSS sg13_hv_nmos W=88.00000000000001 L=0.5999999999999999
* device instance $860 r0 *1 90.95,785.52 sg13_hv_nmos
M$860 VSS \$1282 IN3 VSS sg13_hv_nmos W=88.00000000000001 L=0.5999999999999999
* device instance $880 r0 *1 1209.05,794.58 sg13_hv_nmos
M$880 VSS \$1308 OUT3 VSS sg13_hv_nmos W=35.199999999999996 L=0.5999999999999999
* device instance $888 r0 *1 1064.68,797.64 sg13_hv_nmos
M$888 \$1293 \$1010 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $889 r0 *1 1064.68,798.47 sg13_hv_nmos
M$889 VSS \$1292 \$1302 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $890 r0 *1 1064.68,799.81 sg13_hv_nmos
M$890 VSS \$1302 \$1308 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $891 r0 *1 1064.68,801.15 sg13_hv_nmos
M$891 \$1320 \$1010 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $892 r0 *1 1064.68,801.98 sg13_hv_nmos
M$892 VSS \$1319 \$1327 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $893 r0 *1 1064.68,803.32 sg13_hv_nmos
M$893 VSS \$1327 \$1272 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $894 r0 *1 510.665,859.567 sg13_hv_nmos
M$894 \$1573 \$1573 VSS VSS sg13_hv_nmos W=33.0 L=0.9
* device instance $902 r0 *1 530.16,859.567 sg13_hv_nmos
M$902 \$1575 \$1573 VSS VSS sg13_hv_nmos W=33.0 L=0.9
* device instance $910 r0 *1 495.305,859.662 sg13_hv_nmos
M$910 \$1574 \$1573 VSS VSS sg13_hv_nmos W=33.0 L=0.9
* device instance $918 r0 *1 506.045,858.145 sg13_hv_nmos
M$918 VSS \$1574 \$1648 VSS sg13_hv_nmos W=1.0 L=0.44999999999999996
* device instance $919 r0 *1 495.305,870.8 sg13_hv_nmos
M$919 \$1621 \$1573 \$1648 VSS sg13_hv_nmos W=178.00000000000006
+ L=0.8999999999999999
* device instance $939 r0 *1 540.27,863.82 sg13_hv_nmos
M$939 \$1377 \$1718 \$1575 VSS sg13_hv_nmos W=136.5 L=0.9
* device instance $953 r0 *1 90.95,885.52 sg13_hv_nmos
M$953 VSS \$1736 IN2 VSS sg13_hv_nmos W=88.00000000000001 L=0.5999999999999999
* device instance $973 r0 *1 529.04,863.82 sg13_hv_nmos
M$973 \$1589 VLDO \$1575 VSS sg13_hv_nmos W=136.5 L=0.9
* device instance $987 r0 *1 1064.68,897.64 sg13_hv_nmos
M$987 \$1803 \$1499 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $988 r0 *1 1064.68,898.47 sg13_hv_nmos
M$988 VSS \$1802 \$1812 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $989 r0 *1 1209.05,894.58 sg13_hv_nmos
M$989 VSS \$1818 OUT2 VSS sg13_hv_nmos W=35.199999999999996 L=0.5999999999999999
* device instance $997 r0 *1 1064.68,899.81 sg13_hv_nmos
M$997 VSS \$1812 \$1818 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $998 r0 *1 1064.68,901.15 sg13_hv_nmos
M$998 \$1830 \$1499 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $999 r0 *1 1064.68,901.98 sg13_hv_nmos
M$999 VSS \$1829 \$1837 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1000 r0 *1 1064.68,903.32 sg13_hv_nmos
M$1000 VSS \$1837 \$1712 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1001 r0 *1 90.95,985.52 sg13_hv_nmos
M$1001 VSS \$1906 IN1 VSS sg13_hv_nmos W=88.00000000000001 L=0.5999999999999999
* device instance $1021 r0 *1 1209.05,994.58 sg13_hv_nmos
M$1021 VSS \$1933 OUT1 VSS sg13_hv_nmos W=35.199999999999996
+ L=0.5999999999999999
* device instance $1029 r0 *1 1064.68,997.64 sg13_hv_nmos
M$1029 \$1917 \$1924 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1030 r0 *1 1064.68,998.47 sg13_hv_nmos
M$1030 VSS \$1916 \$1927 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1031 r0 *1 1064.68,999.81 sg13_hv_nmos
M$1031 VSS \$1927 \$1933 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1032 r0 *1 1064.68,1001.15 sg13_hv_nmos
M$1032 \$1945 \$1924 VSS VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1033 r0 *1 1064.68,1001.98 sg13_hv_nmos
M$1033 VSS \$1944 \$1952 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1034 r0 *1 1064.68,1003.32 sg13_hv_nmos
M$1034 VSS \$1952 \$1897 VSS sg13_hv_nmos W=1.9000000000000001
+ L=0.44999999999999996
* device instance $1035 r0 *1 701.765,1060.945 sg13_hv_nmos
M$1035 VSS \$2013 \$2010 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $1036 r0 *1 801.765,1060.945 sg13_hv_nmos
M$1036 VSS \$2014 \$2011 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $1037 r0 *1 901.765,1060.945 sg13_hv_nmos
M$1037 VSS \$2015 \$2012 VSS sg13_hv_nmos W=2.65 L=0.44999999999999996
* device instance $1038 r0 *1 263.22,1139.21 sg13_hv_nmos
M$1038 VSS \$2148 \$2089 VSS sg13_hv_nmos W=108.0 L=0.5
* device instance $1044 r0 *1 273,1139.21 sg13_hv_nmos
M$1044 VSS \$2148 VSS VSS sg13_hv_nmos W=126.0 L=9.5
* device instance $1051 r0 *1 563.22,1139.21 sg13_hv_nmos
M$1051 VSS \$2149 \$2090 VSS sg13_hv_nmos W=108.0 L=0.5
* device instance $1057 r0 *1 573,1139.21 sg13_hv_nmos
M$1057 VSS \$2149 VSS VSS sg13_hv_nmos W=126.0 L=9.5
* device instance $1064 r0 *1 963.22,1139.21 sg13_hv_nmos
M$1064 VSS \$2150 \$2091 VSS sg13_hv_nmos W=108.0 L=0.5
* device instance $1070 r0 *1 973,1139.21 sg13_hv_nmos
M$1070 VSS \$2150 VSS VSS sg13_hv_nmos W=126.0 L=9.5
* device instance $1116 r0 *1 268.155,1194.53 sg13_hv_nmos
M$1116 VSS \$2089 AVDD VSS sg13_hv_nmos W=756.7999999999977 L=0.5999999999999999
* device instance $1159 r0 *1 568.155,1194.53 sg13_hv_nmos
M$1159 VSS \$2090 IOVDD VSS sg13_hv_nmos W=756.7999999999977
+ L=0.5999999999999999
* device instance $1202 r0 *1 968.155,1194.53 sg13_hv_nmos
M$1202 VSS \$2091 VDD VSS sg13_hv_nmos W=756.7999999999977 L=0.5999999999999999
* device instance $1546 r0 *1 385.52,1209.05 sg13_hv_nmos
M$1546 VSS \$2220 VREF VSS sg13_hv_nmos W=88.00000000000001 L=0.5999999999999999
* device instance $1566 r0 *1 485.52,1209.05 sg13_hv_nmos
M$1566 VSS \$2221 VLDO VSS sg13_hv_nmos W=88.00000000000001 L=0.5999999999999999
* device instance $1672 r0 *1 500.255,243.995 sg13_lv_pmos
M$1672 \$181 \$186 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $1673 r0 *1 700.255,243.995 sg13_lv_pmos
M$1673 \$182 \$187 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $1674 r0 *1 800.255,243.995 sg13_lv_pmos
M$1674 \$183 \$188 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $1675 r0 *1 900.255,243.995 sg13_lv_pmos
M$1675 \$184 \$189 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $1676 r0 *1 1056.005,297.48 sg13_lv_pmos
M$1676 \$235 \$237 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $1677 r0 *1 1056.005,300.99 sg13_lv_pmos
M$1677 \$263 \$237 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $1678 r0 *1 1056.005,397.48 sg13_lv_pmos
M$1678 \$350 \$352 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $1679 r0 *1 1056.005,400.99 sg13_lv_pmos
M$1679 \$378 \$352 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $1680 r0 *1 1056.005,497.48 sg13_lv_pmos
M$1680 \$465 \$467 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $1681 r0 *1 1056.005,500.99 sg13_lv_pmos
M$1681 \$493 \$467 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $1682 r0 *1 484.613,506.087 sg13_lv_pmos
M$1682 VDD \$515 \$516 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $1683 r0 *1 485.123,506.087 sg13_lv_pmos
M$1683 \$516 \$527 \$517 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $1684 r0 *1 485.773,506.417 sg13_lv_pmos
M$1684 \$517 \$510 \$551 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1685 r0 *1 486.108,506.417 sg13_lv_pmos
M$1685 \$551 \$518 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1686 r0 *1 486.618,506.417 sg13_lv_pmos
M$1686 VDD \$504 \$518 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1687 r0 *1 487.128,506.417 sg13_lv_pmos
M$1687 VDD \$517 \$518 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1688 r0 *1 487.688,506.252 sg13_lv_pmos
M$1688 VDD \$517 \$519 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1689 r0 *1 497.628,506.266 sg13_lv_pmos
M$1689 VDD \$584 \$534 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $1690 r0 *1 496.608,506.251 sg13_lv_pmos
M$1690 VDD \$534 \$522 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1692 r0 *1 489.163,506.392 sg13_lv_pmos
M$1692 VDD \$517 \$520 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $1693 r0 *1 489.673,506.252 sg13_lv_pmos
M$1693 VDD \$520 \$521 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1694 r0 *1 491.888,506.252 sg13_lv_pmos
M$1694 VDD \$521 \$467 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1696 r0 *1 476.778,506.267 sg13_lv_pmos
M$1696 VDD \$689 \$513 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1697 r0 *1 480.303,506.312 sg13_lv_pmos
M$1697 \$527 \$689 VDD VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $1698 r0 *1 480.813,506.312 sg13_lv_pmos
M$1698 VDD \$527 \$510 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $1699 r0 *1 481.973,506.377 sg13_lv_pmos
M$1699 \$514 \$510 \$515 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1700 r0 *1 482.483,506.377 sg13_lv_pmos
M$1700 \$515 \$527 \$549 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1701 r0 *1 482.858,506.377 sg13_lv_pmos
M$1701 \$549 \$516 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1702 r0 *1 483.433,506.377 sg13_lv_pmos
M$1702 VDD \$504 \$515 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1703 r0 *1 494.703,506.266 sg13_lv_pmos
M$1703 VDD \$181 \$504 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1704 r0 *1 478.773,506.602 sg13_lv_pmos
M$1704 VDD \$584 \$514 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1705 r0 *1 479.283,506.602 sg13_lv_pmos
M$1705 \$514 \$504 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1706 r0 *1 481.401,518.61 sg13_lv_pmos
M$1706 \$581 \$631 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $1707 r0 *1 482.801,518.61 sg13_lv_pmos
M$1707 AVDD \$600 \$581 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $1708 r0 *1 484.201,518.61 sg13_lv_pmos
M$1708 \$600 \$581 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $1709 r0 *1 485.601,518.61 sg13_lv_pmos
M$1709 AVDD \$631 \$600 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $1710 r0 *1 489.122,508.991 sg13_lv_pmos
M$1710 \$564 \$513 \$565 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $1713 r0 *1 488.259,518.61 sg13_lv_pmos
M$1713 \$609 \$600 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $1714 r0 *1 489.659,518.61 sg13_lv_pmos
M$1714 VDD \$584 \$609 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $1715 r0 *1 491.059,518.61 sg13_lv_pmos
M$1715 \$584 \$609 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $1716 r0 *1 492.459,518.61 sg13_lv_pmos
M$1716 VDD \$581 \$584 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $1717 r0 *1 435.35,517.186 sg13_lv_pmos
M$1717 VDD \$686 \$622 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1719 r0 *1 436.38,517.186 sg13_lv_pmos
M$1719 VDD \$633 \$622 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1721 r0 *1 438.155,517.186 sg13_lv_pmos
M$1721 VDD \$622 \$623 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1725 r0 *1 441.035,517.186 sg13_lv_pmos
M$1725 VDD \$623 \$624 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1729 r0 *1 443.915,517.186 sg13_lv_pmos
M$1729 VDD \$624 \$625 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1733 r0 *1 446.795,517.186 sg13_lv_pmos
M$1733 VDD \$625 \$626 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1737 r0 *1 449.675,517.186 sg13_lv_pmos
M$1737 VDD \$626 \$627 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1741 r0 *1 452.555,517.186 sg13_lv_pmos
M$1741 VDD \$627 \$628 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1745 r0 *1 455.51,517.186 sg13_lv_pmos
M$1745 VDD \$628 \$629 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1747 r0 *1 456.54,517.186 sg13_lv_pmos
M$1747 VDD \$626 \$629 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1749 r0 *1 458.315,517.186 sg13_lv_pmos
M$1749 VDD \$629 \$630 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1753 r0 *1 461.135,517.186 sg13_lv_pmos
M$1753 VDD \$630 \$631 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $1761 r0 *1 431.445,522.941 sg13_lv_pmos
M$1761 VDD \$182 \$633 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1763 r0 *1 432.935,536.781 sg13_lv_pmos
M$1763 \$732 \$521 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $1764 r0 *1 433.475,536.921 sg13_lv_pmos
M$1764 VDD \$631 \$733 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1765 r0 *1 433.985,536.921 sg13_lv_pmos
M$1765 \$733 \$732 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1766 r0 *1 433.365,522.941 sg13_lv_pmos
M$1766 VDD \$633 \$679 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1768 r0 *1 435.35,522.941 sg13_lv_pmos
M$1768 VDD \$628 \$707 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1770 r0 *1 436.38,522.941 sg13_lv_pmos
M$1770 VDD \$679 \$707 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1772 r0 *1 438.155,522.941 sg13_lv_pmos
M$1772 VDD \$707 \$681 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1776 r0 *1 441.035,522.941 sg13_lv_pmos
M$1776 VDD \$681 \$682 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1780 r0 *1 443.915,522.941 sg13_lv_pmos
M$1780 VDD \$682 \$683 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1784 r0 *1 446.795,522.941 sg13_lv_pmos
M$1784 VDD \$683 \$684 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1788 r0 *1 449.675,522.941 sg13_lv_pmos
M$1788 VDD \$684 \$685 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1792 r0 *1 452.555,522.941 sg13_lv_pmos
M$1792 VDD \$685 \$686 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1796 r0 *1 455.51,522.941 sg13_lv_pmos
M$1796 VDD \$686 \$692 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1798 r0 *1 456.54,522.941 sg13_lv_pmos
M$1798 VDD \$684 \$692 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1800 r0 *1 458.315,522.941 sg13_lv_pmos
M$1800 VDD \$692 \$688 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1804 r0 *1 461.135,522.941 sg13_lv_pmos
M$1804 VDD \$688 \$689 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $1812 r0 *1 467.935,536.781 sg13_lv_pmos
M$1812 \$738 \$522 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $1813 r0 *1 468.475,536.921 sg13_lv_pmos
M$1813 VDD \$689 \$739 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1814 r0 *1 468.985,536.921 sg13_lv_pmos
M$1814 \$739 \$738 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1815 r0 *1 431.51,536.936 sg13_lv_pmos
M$1815 VDD \$689 \$731 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1816 r0 *1 435.785,537.061 sg13_lv_pmos
M$1816 VDD \$631 \$734 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $1817 r0 *1 436.295,537.061 sg13_lv_pmos
M$1817 VDD \$521 \$734 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $1818 r0 *1 436.805,536.921 sg13_lv_pmos
M$1818 VDD \$734 \$735 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1819 r0 *1 452.577,539.206 sg13_lv_pmos
M$1819 \$752 \$757 AVDD AVDD sg13_lv_pmos W=10.5 L=1.5
* device instance $1823 r0 *1 466.51,536.936 sg13_lv_pmos
M$1823 VDD \$631 \$737 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1824 r0 *1 470.785,537.061 sg13_lv_pmos
M$1824 VDD \$689 \$740 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $1825 r0 *1 471.295,537.061 sg13_lv_pmos
M$1825 VDD \$522 \$740 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $1826 r0 *1 471.805,536.921 sg13_lv_pmos
M$1826 VDD \$740 \$741 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1827 r0 *1 487.577,539.206 sg13_lv_pmos
M$1827 \$564 \$758 AVDD AVDD sg13_lv_pmos W=10.5 L=1.5
* device instance $1831 r0 *1 440.927,539.221 sg13_lv_pmos
M$1831 \$736 \$736 AVDD AVDD sg13_lv_pmos W=10.5 L=1.5
* device instance $1835 r0 *1 475.927,539.221 sg13_lv_pmos
M$1835 \$569 \$569 AVDD AVDD sg13_lv_pmos W=10.5 L=1.5
* device instance $1839 r0 *1 434.41,549.416 sg13_lv_pmos
M$1839 \$791 \$733 VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $1840 r0 *1 436.765,548.916 sg13_lv_pmos
M$1840 \$791 \$731 \$587 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $1843 r0 *1 469.41,549.416 sg13_lv_pmos
M$1843 \$792 \$739 VHI AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $1844 r0 *1 471.765,548.916 sg13_lv_pmos
M$1844 \$792 \$737 \$752 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $1847 r0 *1 449.83,598.84 sg13_lv_pmos
M$1847 VDD \$910 \$868 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1849 r0 *1 450.86,598.84 sg13_lv_pmos
M$1849 VDD \$867 \$868 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1851 r0 *1 452.635,598.84 sg13_lv_pmos
M$1851 VDD \$868 \$858 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1855 r0 *1 455.515,598.84 sg13_lv_pmos
M$1855 VDD \$858 \$859 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1859 r0 *1 458.395,598.84 sg13_lv_pmos
M$1859 VDD \$859 \$860 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1863 r0 *1 461.275,598.84 sg13_lv_pmos
M$1863 VDD \$860 \$861 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1867 r0 *1 464.155,598.84 sg13_lv_pmos
M$1867 VDD \$861 \$862 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1871 r0 *1 467.035,598.84 sg13_lv_pmos
M$1871 VDD \$862 \$863 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1875 r0 *1 469.99,598.84 sg13_lv_pmos
M$1875 VDD \$863 \$869 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1877 r0 *1 471.02,598.84 sg13_lv_pmos
M$1877 VDD \$861 \$869 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1879 r0 *1 472.795,598.84 sg13_lv_pmos
M$1879 VDD \$869 \$865 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1883 r0 *1 475.615,598.84 sg13_lv_pmos
M$1883 VDD \$865 \$866 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $1891 r0 *1 445.925,604.64 sg13_lv_pmos
M$1891 VDD \$853 \$867 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1893 r0 *1 447.845,604.64 sg13_lv_pmos
M$1893 VDD \$867 \$903 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1895 r0 *1 449.83,604.64 sg13_lv_pmos
M$1895 VDD \$863 \$914 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1897 r0 *1 450.86,604.64 sg13_lv_pmos
M$1897 VDD \$903 \$914 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1899 r0 *1 452.635,604.64 sg13_lv_pmos
M$1899 VDD \$914 \$905 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1903 r0 *1 455.515,604.64 sg13_lv_pmos
M$1903 VDD \$905 \$906 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1907 r0 *1 458.395,604.64 sg13_lv_pmos
M$1907 VDD \$906 \$907 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1911 r0 *1 461.275,604.64 sg13_lv_pmos
M$1911 VDD \$907 \$908 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1915 r0 *1 464.155,604.64 sg13_lv_pmos
M$1915 VDD \$908 \$909 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1919 r0 *1 467.035,604.64 sg13_lv_pmos
M$1919 VDD \$909 \$910 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1923 r0 *1 469.99,604.64 sg13_lv_pmos
M$1923 VDD \$910 \$915 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1925 r0 *1 471.02,604.64 sg13_lv_pmos
M$1925 VDD \$908 \$915 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1927 r0 *1 472.795,604.64 sg13_lv_pmos
M$1927 VDD \$915 \$912 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $1931 r0 *1 475.615,604.64 sg13_lv_pmos
M$1931 VDD \$912 \$913 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $1939 r0 *1 433.28,618.09 sg13_lv_pmos
M$1939 VDD \$913 \$975 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1940 r0 *1 434.36,617.935 sg13_lv_pmos
M$1940 \$979 \$946 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $1941 r0 *1 434.9,618.075 sg13_lv_pmos
M$1941 VDD \$866 \$976 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1942 r0 *1 435.41,618.075 sg13_lv_pmos
M$1942 \$976 \$979 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1943 r0 *1 434.995,621.675 sg13_lv_pmos
M$1943 \$1344 \$975 \$1015 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $1946 r0 *1 436.85,618.215 sg13_lv_pmos
M$1946 VDD \$866 \$984 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $1947 r0 *1 437.36,618.215 sg13_lv_pmos
M$1947 VDD \$946 \$984 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $1948 r0 *1 437.87,618.075 sg13_lv_pmos
M$1948 VDD \$984 \$967 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1949 r0 *1 439.97,617.765 sg13_lv_pmos
M$1949 VHI \$976 \$1015 AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $1950 r0 *1 469.335,618.09 sg13_lv_pmos
M$1950 VDD \$866 \$977 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1951 r0 *1 470.415,617.935 sg13_lv_pmos
M$1951 \$980 \$947 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $1952 r0 *1 470.955,618.075 sg13_lv_pmos
M$1952 VDD \$913 \$978 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1953 r0 *1 471.465,618.075 sg13_lv_pmos
M$1953 \$978 \$980 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1954 r0 *1 471.05,621.675 sg13_lv_pmos
M$1954 \$1016 \$977 \$1017 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $1957 r0 *1 472.905,618.215 sg13_lv_pmos
M$1957 VDD \$913 \$985 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $1958 r0 *1 473.415,618.215 sg13_lv_pmos
M$1958 VDD \$947 \$985 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $1959 r0 *1 473.925,618.075 sg13_lv_pmos
M$1959 VDD \$985 \$969 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1960 r0 *1 476.025,617.765 sg13_lv_pmos
M$1960 VHI \$978 \$1017 AVDD sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $1961 r0 *1 505.435,618.205 sg13_lv_pmos
M$1961 VDD \$913 \$981 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1962 r0 *1 520.805,621.42 sg13_lv_pmos
M$1962 VDD \$1047 \$1037 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1963 r0 *1 521.315,621.42 sg13_lv_pmos
M$1963 VDD \$1033 \$1037 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1964 r0 *1 521.765,621.71 sg13_lv_pmos
M$1964 VDD \$1062 \$1038 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $1965 r0 *1 526.15,621.66 sg13_lv_pmos
M$1965 \$1073 \$1039 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1966 r0 *1 526.875,621.66 sg13_lv_pmos
M$1966 VDD \$913 \$1039 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1967 r0 *1 529.005,621.405 sg13_lv_pmos
M$1967 \$1048 \$1073 \$1084 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1968 r0 *1 529.385,621.405 sg13_lv_pmos
M$1968 \$1084 \$1041 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1969 r0 *1 529.995,621.405 sg13_lv_pmos
M$1969 VDD \$1033 \$1041 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1970 r0 *1 530.505,621.405 sg13_lv_pmos
M$1970 VDD \$1048 \$1041 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $1971 r0 *1 532.065,621.51 sg13_lv_pmos
M$1971 VDD \$1048 \$1043 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $1972 r0 *1 531.045,621.57 sg13_lv_pmos
M$1972 VDD \$1048 \$1042 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1974 r0 *1 528.31,621.695 sg13_lv_pmos
M$1974 \$1038 \$1039 \$1048 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $1975 r0 *1 533.15,621.67 sg13_lv_pmos
M$1975 VDD \$1043 \$946 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1977 r0 *1 535.2,621.67 sg13_lv_pmos
M$1977 VDD \$946 \$1010 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $1979 r0 *1 536.99,621.68 sg13_lv_pmos
M$1979 \$1033 \$181 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $1980 r0 *1 456.64,625.975 sg13_lv_pmos
M$1980 \$1016 \$1105 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $1984 r0 *1 462.64,625.975 sg13_lv_pmos
M$1984 \$968 \$968 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $1988 r0 *1 492.695,625.975 sg13_lv_pmos
M$1988 \$1018 \$1106 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $1992 r0 *1 498.695,625.975 sg13_lv_pmos
M$1992 \$970 \$970 AVDD AVDD sg13_lv_pmos W=10.0 L=1.5
* device instance $1996 r0 *1 505.15,621.115 sg13_lv_pmos
M$1996 \$1061 \$981 \$1018 AVDD sg13_lv_pmos W=6.0 L=0.13
* device instance $1999 r0 *1 521.51,632.615 sg13_lv_pmos
M$1999 VDD \$1134 \$1129 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2000 r0 *1 522.815,621.785 sg13_lv_pmos
M$2000 \$1062 \$1033 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2001 r0 *1 523.55,621.785 sg13_lv_pmos
M$2001 VDD \$1038 \$1083 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2002 r0 *1 523.94,621.785 sg13_lv_pmos
M$2002 \$1083 \$1039 \$1062 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2003 r0 *1 524.45,621.785 sg13_lv_pmos
M$2003 \$1062 \$1073 \$1037 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2004 r0 *1 524.18,632.615 sg13_lv_pmos
M$2004 \$1129 \$1047 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2005 r0 *1 528.19,632.615 sg13_lv_pmos
M$2005 VDD \$1129 \$1047 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2006 r0 *1 530.86,632.615 sg13_lv_pmos
M$2006 \$1047 \$1133 VDD VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2007 r0 *1 534.455,625.47 sg13_lv_pmos
M$2007 VDD \$1103 \$947 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2009 r0 *1 534.47,626.49 sg13_lv_pmos
M$2009 VDD \$1047 \$1103 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2010 r0 *1 508.41,633.315 sg13_lv_pmos
M$2010 AVDD \$866 \$1133 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2011 r0 *1 511.055,633.315 sg13_lv_pmos
M$2011 \$1133 \$1134 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2012 r0 *1 513.41,633.315 sg13_lv_pmos
M$2012 AVDD \$1133 \$1134 AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2013 r0 *1 516.045,633.315 sg13_lv_pmos
M$2013 \$1134 \$866 AVDD AVDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2014 r0 *1 1056.005,797.48 sg13_lv_pmos
M$2014 \$1292 \$1010 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2015 r0 *1 1056.005,800.99 sg13_lv_pmos
M$2015 \$1319 \$1010 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2016 r0 *1 633.21,840.21 sg13_lv_pmos
M$2016 VLDO \$1380 \$1380 VLDO sg13_lv_pmos W=10.0 L=1.5
* device instance $2018 r0 *1 630.06,845.38 sg13_lv_pmos
M$2018 \$1391 \$1422 \$1384 VLDO sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2020 r0 *1 622.075,848.775 sg13_lv_pmos
M$2020 VLDO \$1457 \$1413 VLDO sg13_lv_pmos W=4.0 L=0.13
* device instance $2022 r0 *1 624.015,848.775 sg13_lv_pmos
M$2022 VLDO \$1412 \$1413 VLDO sg13_lv_pmos W=4.0 L=0.13
* device instance $2024 r0 *1 625.955,848.775 sg13_lv_pmos
M$2024 VLDO \$1413 \$1412 VLDO sg13_lv_pmos W=4.0 L=0.13
* device instance $2026 r0 *1 627.895,848.775 sg13_lv_pmos
M$2026 VLDO \$1457 \$1412 VLDO sg13_lv_pmos W=4.0 L=0.13
* device instance $2028 r0 *1 631.3,848.775 sg13_lv_pmos
M$2028 VDD \$1412 \$1419 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2030 r0 *1 633.24,848.775 sg13_lv_pmos
M$2030 VDD \$1414 \$1419 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2032 r0 *1 635.18,848.775 sg13_lv_pmos
M$2032 VDD \$1419 \$1414 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2034 r0 *1 637.12,848.775 sg13_lv_pmos
M$2034 VDD \$1413 \$1414 VDD sg13_lv_pmos W=4.0 L=0.13
* device instance $2036 r0 *1 585.345,849.525 sg13_lv_pmos
M$2036 \$1417 \$1473 \$1854 VLDO sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2038 r0 *1 586.14,853.855 sg13_lv_pmos
M$2038 VHI \$1533 \$1417 VLDO sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2039 r0 *1 592.87,850.555 sg13_lv_pmos
M$2039 VLDO \$1386 \$1406 VLDO sg13_lv_pmos W=10.0 L=1.5
* device instance $2041 r0 *1 606.935,849.525 sg13_lv_pmos
M$2041 \$1418 \$1474 \$1406 VLDO sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $2043 r0 *1 607.73,853.855 sg13_lv_pmos
M$2043 VHI \$1534 \$1418 VLDO sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $2044 r0 *1 614.46,850.555 sg13_lv_pmos
M$2044 VLDO \$1387 \$1391 VLDO sg13_lv_pmos W=10.0 L=1.5
* device instance $2046 r0 *1 628.87,853.995 sg13_lv_pmos
M$2046 \$1506 \$1493 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2047 r0 *1 629.595,853.995 sg13_lv_pmos
M$2047 VDD \$1434 \$1493 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2048 r0 *1 620.95,854.02 sg13_lv_pmos
M$2048 VDD \$1434 \$1422 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2049 r0 *1 622.39,854.02 sg13_lv_pmos
M$2049 VDD \$181 \$1489 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2050 r0 *1 635.87,854.005 sg13_lv_pmos
M$2050 VDD \$1497 \$1590 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2052 r0 *1 637.86,854.02 sg13_lv_pmos
M$2052 VDD \$1414 \$1498 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2053 r0 *1 638.37,854.005 sg13_lv_pmos
M$2053 VDD \$1498 \$1591 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2055 r0 *1 640.39,854.005 sg13_lv_pmos
M$2055 VDD \$1590 \$1499 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2057 r0 *1 617.465,865.11 sg13_lv_pmos
M$2057 VDD \$1626 \$1607 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2059 r0 *1 618.495,865.11 sg13_lv_pmos
M$2059 VDD \$1627 \$1607 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2061 r0 *1 623.525,853.755 sg13_lv_pmos
M$2061 VDD \$1414 \$1490 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2062 r0 *1 624.035,853.755 sg13_lv_pmos
M$2062 VDD \$1489 \$1490 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2063 r0 *1 624.485,854.045 sg13_lv_pmos
M$2063 VDD \$1535 \$1491 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2064 r0 *1 625.535,854.12 sg13_lv_pmos
M$2064 \$1535 \$1489 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2065 r0 *1 626.27,854.12 sg13_lv_pmos
M$2065 VDD \$1491 \$1554 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2066 r0 *1 626.66,854.12 sg13_lv_pmos
M$2066 \$1554 \$1493 \$1535 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2067 r0 *1 627.17,854.12 sg13_lv_pmos
M$2067 \$1535 \$1506 \$1490 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2068 r0 *1 631.725,853.74 sg13_lv_pmos
M$2068 \$1507 \$1506 \$1549 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2069 r0 *1 632.105,853.74 sg13_lv_pmos
M$2069 \$1549 \$1495 VDD VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2070 r0 *1 632.715,853.74 sg13_lv_pmos
M$2070 VDD \$1489 \$1495 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2071 r0 *1 633.225,853.74 sg13_lv_pmos
M$2071 VDD \$1507 \$1495 VDD sg13_lv_pmos W=0.42 L=0.13
* device instance $2072 r0 *1 634.785,853.845 sg13_lv_pmos
M$2072 VDD \$1507 \$1497 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2073 r0 *1 633.765,853.905 sg13_lv_pmos
M$2073 VDD \$1507 \$1496 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2075 r0 *1 631.03,854.03 sg13_lv_pmos
M$2075 \$1491 \$1493 \$1507 VDD sg13_lv_pmos W=1.0 L=0.13
* device instance $2076 r0 *1 640.7,865.11 sg13_lv_pmos
M$2076 VDD \$1597 \$1608 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2078 r0 *1 641.73,865.11 sg13_lv_pmos
M$2078 VDD \$1596 \$1608 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2080 r0 *1 643.75,865.11 sg13_lv_pmos
M$2080 VDD \$1608 \$1599 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2084 r0 *1 623.374,865.112 sg13_lv_pmos
M$2084 VDD \$1593 \$1594 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2088 r0 *1 626.254,865.112 sg13_lv_pmos
M$2088 VDD \$1594 \$1595 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2092 r0 *1 629.134,865.112 sg13_lv_pmos
M$2092 VDD \$1595 \$1596 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2096 r0 *1 632.714,865.112 sg13_lv_pmos
M$2096 VDD \$1596 \$1458 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2100 r0 *1 636.294,865.112 sg13_lv_pmos
M$2100 VDD \$1458 \$1597 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2104 r0 *1 646.57,865.112 sg13_lv_pmos
M$2104 VDD \$1599 \$1457 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2112 r0 *1 577.495,865.995 sg13_lv_pmos
M$2112 VDD \$1457 \$1622 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2113 r0 *1 578.005,865.995 sg13_lv_pmos
M$2113 VDD \$1590 \$1622 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2114 r0 *1 578.515,865.855 sg13_lv_pmos
M$2114 VDD \$1622 \$1504 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2115 r0 *1 579.805,865.715 sg13_lv_pmos
M$2115 \$1623 \$1590 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2116 r0 *1 580.345,865.855 sg13_lv_pmos
M$2116 VDD \$1457 \$1533 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2117 r0 *1 580.855,865.855 sg13_lv_pmos
M$2117 \$1533 \$1623 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2118 r0 *1 582.565,865.87 sg13_lv_pmos
M$2118 VDD \$1434 \$1473 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2119 r0 *1 599.085,865.995 sg13_lv_pmos
M$2119 VDD \$1434 \$1624 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2120 r0 *1 599.595,865.995 sg13_lv_pmos
M$2120 VDD \$1591 \$1624 VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2121 r0 *1 600.105,865.855 sg13_lv_pmos
M$2121 VDD \$1624 \$1505 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2122 r0 *1 601.395,865.715 sg13_lv_pmos
M$2122 \$1625 \$1591 VDD VDD sg13_lv_pmos W=0.84 L=0.13
* device instance $2123 r0 *1 601.935,865.855 sg13_lv_pmos
M$2123 VDD \$1434 \$1534 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2124 r0 *1 602.445,865.855 sg13_lv_pmos
M$2124 \$1534 \$1625 VDD VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2125 r0 *1 604.155,865.87 sg13_lv_pmos
M$2125 VDD \$1457 \$1474 VDD sg13_lv_pmos W=1.12 L=0.13
* device instance $2126 r0 *1 620.494,870.782 sg13_lv_pmos
M$2126 VDD \$1678 \$1671 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2130 r0 *1 620.494,865.114 sg13_lv_pmos
M$2130 VDD \$1607 \$1593 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2134 r0 *1 623.374,870.782 sg13_lv_pmos
M$2134 VDD \$1671 \$1672 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2138 r0 *1 626.254,870.782 sg13_lv_pmos
M$2138 VDD \$1672 \$1673 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2142 r0 *1 629.134,870.782 sg13_lv_pmos
M$2142 VDD \$1673 \$1674 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2146 r0 *1 632.714,870.782 sg13_lv_pmos
M$2146 VDD \$1674 \$1675 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2150 r0 *1 636.294,870.782 sg13_lv_pmos
M$2150 VDD \$1675 \$1626 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2154 r0 *1 643.505,870.782 sg13_lv_pmos
M$2154 VDD \$1679 \$1677 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $2158 r0 *1 613.56,870.787 sg13_lv_pmos
M$2158 VDD \$1692 \$1627 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2160 r0 *1 615.48,870.787 sg13_lv_pmos
M$2160 VDD \$1627 \$1669 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2162 r0 *1 617.465,870.787 sg13_lv_pmos
M$2162 VDD \$1597 \$1678 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2164 r0 *1 618.495,870.787 sg13_lv_pmos
M$2164 VDD \$1669 \$1678 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2166 r0 *1 640.44,870.787 sg13_lv_pmos
M$2166 VDD \$1626 \$1679 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2168 r0 *1 641.47,870.787 sg13_lv_pmos
M$2168 VDD \$1674 \$1679 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $2170 r0 *1 646.325,870.788 sg13_lv_pmos
M$2170 VDD \$1677 \$1434 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $2178 r0 *1 1056.005,897.48 sg13_lv_pmos
M$2178 \$1802 \$1499 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2179 r0 *1 1056.005,900.99 sg13_lv_pmos
M$2179 \$1829 \$1499 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2180 r0 *1 1056.005,997.48 sg13_lv_pmos
M$2180 \$1916 \$1924 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2181 r0 *1 1056.005,1000.99 sg13_lv_pmos
M$2181 \$1944 \$1924 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2182 r0 *1 700.255,1056.005 sg13_lv_pmos
M$2182 \$853 \$2010 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2183 r0 *1 800.255,1056.005 sg13_lv_pmos
M$2183 \$1692 \$2011 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2184 r0 *1 900.255,1056.005 sg13_lv_pmos
M$2184 \$2005 \$2012 VDD VDD sg13_lv_pmos W=4.75 L=0.12999999999999998
* device instance $2185 r0 *1 501.765,243.945 sg13_hv_pmos
M$2185 VDD \$129 \$186 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $2186 r0 *1 701.765,243.945 sg13_hv_pmos
M$2186 VDD \$130 \$187 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $2187 r0 *1 801.765,243.945 sg13_hv_pmos
M$2187 VDD \$132 \$188 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $2188 r0 *1 901.765,243.945 sg13_hv_pmos
M$2188 VDD \$133 \$189 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $2189 r0 *1 151.08,285.52 sg13_hv_pmos
M$2189 AVDD \$226 IN6 AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $2229 r0 *1 1141.82,294.58 sg13_hv_pmos
M$2229 IOVDD \$216 OUT6 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $2245 r0 *1 1068.82,297.64 sg13_hv_pmos
M$2245 \$236 \$246 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2246 r0 *1 1068.82,298.47 sg13_hv_pmos
M$2246 IOVDD \$236 \$246 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2247 r0 *1 1068.82,299.81 sg13_hv_pmos
M$2247 IOVDD \$246 \$252 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $2248 r0 *1 1068.82,301.15 sg13_hv_pmos
M$2248 \$264 \$271 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2249 r0 *1 1068.82,301.98 sg13_hv_pmos
M$2249 IOVDD \$264 \$271 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2250 r0 *1 1068.82,303.32 sg13_hv_pmos
M$2250 IOVDD \$271 \$216 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $2251 r0 *1 151.08,385.52 sg13_hv_pmos
M$2251 AVDD \$341 IN5 AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $2291 r0 *1 1141.82,394.58 sg13_hv_pmos
M$2291 IOVDD \$331 OUT5 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $2307 r0 *1 1068.82,397.64 sg13_hv_pmos
M$2307 \$351 \$361 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2308 r0 *1 1068.82,398.47 sg13_hv_pmos
M$2308 IOVDD \$351 \$361 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2309 r0 *1 1068.82,399.81 sg13_hv_pmos
M$2309 IOVDD \$361 \$367 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $2310 r0 *1 1068.82,401.15 sg13_hv_pmos
M$2310 \$379 \$386 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2311 r0 *1 1068.82,401.98 sg13_hv_pmos
M$2311 IOVDD \$379 \$386 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2312 r0 *1 1068.82,403.32 sg13_hv_pmos
M$2312 IOVDD \$386 \$331 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $2313 r0 *1 151.08,485.52 sg13_hv_pmos
M$2313 AVDD \$456 IN4 AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $2353 r0 *1 1141.82,494.58 sg13_hv_pmos
M$2353 IOVDD \$446 OUT4 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $2369 r0 *1 1068.82,497.64 sg13_hv_pmos
M$2369 \$466 \$476 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2370 r0 *1 1068.82,498.47 sg13_hv_pmos
M$2370 IOVDD \$466 \$476 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2371 r0 *1 1068.82,499.81 sg13_hv_pmos
M$2371 IOVDD \$476 \$482 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $2372 r0 *1 1068.82,501.15 sg13_hv_pmos
M$2372 \$494 \$501 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2373 r0 *1 1068.82,501.98 sg13_hv_pmos
M$2373 IOVDD \$494 \$501 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2374 r0 *1 1068.82,503.32 sg13_hv_pmos
M$2374 IOVDD \$501 \$446 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $2375 r0 *1 151.08,585.52 sg13_hv_pmos
M$2375 AVDD \$846 VLO AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $2415 r0 *1 151.08,685.52 sg13_hv_pmos
M$2415 AVDD \$1191 VHI AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $2455 r0 *1 1125.09,678.44 sg13_hv_pmos
M$2455 IOVDD \$1185 \$1184 IOVDD sg13_hv_pmos W=350.0 L=0.5
* device instance $2505 r0 *1 151.08,785.52 sg13_hv_pmos
M$2505 AVDD \$1283 IN3 AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $2545 r0 *1 1141.82,794.58 sg13_hv_pmos
M$2545 IOVDD \$1272 OUT3 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $2561 r0 *1 1068.82,797.64 sg13_hv_pmos
M$2561 \$1293 \$1302 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2562 r0 *1 1068.82,798.47 sg13_hv_pmos
M$2562 IOVDD \$1293 \$1302 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2563 r0 *1 1068.82,799.81 sg13_hv_pmos
M$2563 IOVDD \$1302 \$1308 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $2564 r0 *1 1068.82,801.15 sg13_hv_pmos
M$2564 \$1320 \$1327 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2565 r0 *1 1068.82,801.98 sg13_hv_pmos
M$2565 IOVDD \$1320 \$1327 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2566 r0 *1 1068.82,803.32 sg13_hv_pmos
M$2566 IOVDD \$1327 \$1272 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $2567 r0 *1 519.105,828.1 sg13_hv_pmos
M$2567 IOVDD \$1377 VLDO IOVDD sg13_hv_pmos W=1414.0 L=0.44999999999999996
* device instance $2595 r0 *1 497.865,880.705 sg13_hv_pmos
M$2595 IOVDD \$1648 \$1648 IOVDD sg13_hv_pmos W=54.0 L=0.8999999999999999
* device instance $2613 r0 *1 495.265,883.64 sg13_hv_pmos
M$2613 \$1574 \$1574 IOVDD IOVDD sg13_hv_pmos W=1.0 L=5.0
* device instance $2614 r0 *1 497.865,886.92 sg13_hv_pmos
M$2614 IOVDD \$1648 \$1573 IOVDD sg13_hv_pmos W=54.0 L=0.8999999999999999
* device instance $2632 r0 *1 527.575,885.93 sg13_hv_pmos
M$2632 IOVDD \$1589 \$1589 IOVDD sg13_hv_pmos W=36.0 L=0.8999999999999999
* device instance $2638 r0 *1 535.255,885.93 sg13_hv_pmos
M$2638 IOVDD \$1589 \$1377 IOVDD sg13_hv_pmos W=36.0 L=0.8999999999999999
* device instance $2644 r0 *1 151.08,885.52 sg13_hv_pmos
M$2644 AVDD \$1737 IN2 AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $2684 r0 *1 1068.82,899.81 sg13_hv_pmos
M$2684 IOVDD \$1812 \$1818 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $2685 r0 *1 1068.82,897.64 sg13_hv_pmos
M$2685 \$1803 \$1812 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2686 r0 *1 1068.82,898.47 sg13_hv_pmos
M$2686 IOVDD \$1803 \$1812 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2687 r0 *1 1141.82,894.58 sg13_hv_pmos
M$2687 IOVDD \$1712 OUT2 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $2703 r0 *1 1068.82,901.15 sg13_hv_pmos
M$2703 \$1830 \$1837 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2704 r0 *1 1068.82,901.98 sg13_hv_pmos
M$2704 IOVDD \$1830 \$1837 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2705 r0 *1 1068.82,903.32 sg13_hv_pmos
M$2705 IOVDD \$1837 \$1712 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $2706 r0 *1 151.08,985.52 sg13_hv_pmos
M$2706 AVDD \$1907 IN1 AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $2746 r0 *1 1141.82,994.58 sg13_hv_pmos
M$2746 IOVDD \$1897 OUT1 IOVDD sg13_hv_pmos W=106.55999999999996 L=0.6
* device instance $2762 r0 *1 1068.82,997.64 sg13_hv_pmos
M$2762 \$1917 \$1927 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2763 r0 *1 1068.82,998.47 sg13_hv_pmos
M$2763 IOVDD \$1917 \$1927 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2764 r0 *1 1068.82,999.81 sg13_hv_pmos
M$2764 IOVDD \$1927 \$1933 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $2765 r0 *1 1068.82,1001.15 sg13_hv_pmos
M$2765 \$1945 \$1952 IOVDD IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2766 r0 *1 1068.82,1001.98 sg13_hv_pmos
M$2766 IOVDD \$1945 \$1952 IOVDD sg13_hv_pmos W=0.3 L=0.44999999999999996
* device instance $2767 r0 *1 1068.82,1003.32 sg13_hv_pmos
M$2767 IOVDD \$1952 \$1897 IOVDD sg13_hv_pmos W=3.9 L=0.44999999999999996
* device instance $2768 r0 *1 701.765,1056.055 sg13_hv_pmos
M$2768 VDD \$2013 \$2010 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $2769 r0 *1 801.765,1056.055 sg13_hv_pmos
M$2769 VDD \$2014 \$2011 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $2770 r0 *1 901.765,1056.055 sg13_hv_pmos
M$2770 VDD \$2015 \$2012 VDD sg13_hv_pmos W=4.65 L=0.4499999999999999
* device instance $2771 r0 *1 278.44,1125.09 sg13_hv_pmos
M$2771 AVDD \$2148 \$2089 AVDD sg13_hv_pmos W=350.0 L=0.5
* device instance $2821 r0 *1 578.44,1125.09 sg13_hv_pmos
M$2821 IOVDD \$2149 \$2090 IOVDD sg13_hv_pmos W=350.0 L=0.5
* device instance $2871 r0 *1 978.44,1125.09 sg13_hv_pmos
M$2871 IOVDD \$2150 \$2091 IOVDD sg13_hv_pmos W=350.0 L=0.5
* device instance $2921 r0 *1 385.52,1148.92 sg13_hv_pmos
M$2921 AVDD \$2106 VREF AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $2961 r0 *1 485.52,1141.82 sg13_hv_pmos
M$2961 AVDD \$2107 VLDO AVDD sg13_hv_pmos W=266.3999999999999 L=0.6
* device instance $3001 r0 *1 264.54,104.19 dantenna
D$3001 VSS VSS dantenna A=35.0028 P=58.08 m=10
* device instance $3005 r0 *1 464.54,104.19 dantenna
D$3005 VSS RES dantenna A=35.0028 P=58.08 m=2
* device instance $3009 r0 *1 664.54,104.19 dantenna
D$3009 VSS CK4 dantenna A=35.0028 P=58.08 m=2
* device instance $3011 r0 *1 764.54,104.19 dantenna
D$3011 VSS CK5 dantenna A=35.0028 P=58.08 m=2
* device instance $3013 r0 *1 864.54,104.19 dantenna
D$3013 VSS CK6 dantenna A=35.0028 P=58.08 m=2
* device instance $3017 r0 *1 100.44,400 dantenna
D$3017 VSS IN5 dantenna A=35.0028 P=58.08 m=2
* device instance $3018 r0 *1 100.44,300 dantenna
D$3018 VSS IN6 dantenna A=35.0028 P=58.08 m=2
* device instance $3021 r0 *1 222.54,417.63 dantenna
D$3021 VSS \$403 dantenna A=1.984 P=7.48 m=1
* device instance $3022 r0 *1 222.54,317.63 dantenna
D$3022 VSS \$288 dantenna A=1.984 P=7.48 m=1
* device instance $3023 r0 *1 505.225,222.54 dantenna
D$3023 VSS \$129 dantenna A=1.984 P=7.48 m=1
* device instance $3024 r0 *1 705.225,222.54 dantenna
D$3024 VSS \$130 dantenna A=1.984 P=7.48 m=1
* device instance $3025 r0 *1 805.225,222.54 dantenna
D$3025 VSS \$132 dantenna A=1.984 P=7.48 m=1
* device instance $3026 r0 *1 905.225,222.54 dantenna
D$3026 VSS \$133 dantenna A=1.984 P=7.48 m=1
* device instance $3027 r0 *1 1195.06,300 dantenna
D$3027 VSS OUT6 dantenna A=35.0028 P=58.08 m=2
* device instance $3028 r0 *1 1195.06,400 dantenna
D$3028 VSS OUT5 dantenna A=35.0028 P=58.08 m=2
* device instance $3031 r0 *1 1207.17,377.975 dantenna
D$3031 VSS \$367 dantenna A=0.192 P=1.88 m=1
* device instance $3032 r0 *1 1207.17,277.975 dantenna
D$3032 VSS \$252 dantenna A=0.192 P=1.88 m=1
* device instance $3033 r0 *1 1207.17,477.975 dantenna
D$3033 VSS \$482 dantenna A=0.192 P=1.88 m=1
* device instance $3034 r0 *1 100.44,500 dantenna
D$3034 VSS IN4 dantenna A=35.0028 P=58.08 m=2
* device instance $3036 r0 *1 1195.06,500 dantenna
D$3036 VSS OUT4 dantenna A=35.0028 P=58.08 m=2
* device instance $3038 r0 *1 222.54,517.63 dantenna
D$3038 VSS \$587 dantenna A=1.984 P=7.48 m=1
* device instance $3041 r0 *1 100.44,600 dantenna
D$3041 VSS VLO dantenna A=35.0028 P=58.08 m=2
* device instance $3043 r0 *1 222.54,617.63 dantenna
D$3043 VSS \$953 dantenna A=1.984 P=7.48 m=1
* device instance $3044 r0 *1 1192.65,664.765 dantenna
D$3044 VSS \$1184 dantenna A=0.192 P=1.88 m=1
* device instance $3045 r0 *1 100.44,700 dantenna
D$3045 VSS VHI dantenna A=35.0028 P=58.08 m=2
* device instance $3047 r0 *1 222.54,717.63 dantenna
D$3047 VSS \$1218 dantenna A=1.984 P=7.48 m=1
* device instance $3048 r0 *1 1207.17,777.975 dantenna
D$3048 VSS \$1308 dantenna A=0.192 P=1.88 m=1
* device instance $3049 r0 *1 100.44,800 dantenna
D$3049 VSS IN3 dantenna A=35.0028 P=58.08 m=2
* device instance $3051 r0 *1 1195.06,800 dantenna
D$3051 VSS OUT3 dantenna A=35.0028 P=58.08 m=2
* device instance $3053 r0 *1 222.54,817.63 dantenna
D$3053 VSS \$1344 dantenna A=1.984 P=7.48 m=1
* device instance $3054 r0 *1 1207.17,877.975 dantenna
D$3054 VSS \$1818 dantenna A=0.192 P=1.88 m=1
* device instance $3055 r0 *1 100.44,900 dantenna
D$3055 VSS IN2 dantenna A=35.0028 P=58.08 m=2
* device instance $3057 r0 *1 1195.06,900 dantenna
D$3057 VSS OUT2 dantenna A=35.0028 P=58.08 m=2
* device instance $3059 r0 *1 222.54,917.63 dantenna
D$3059 VSS \$1854 dantenna A=1.984 P=7.48 m=1
* device instance $3060 r0 *1 1207.17,977.975 dantenna
D$3060 VSS \$1933 dantenna A=0.192 P=1.88 m=1
* device instance $3061 r0 *1 100.44,1000 dantenna
D$3061 VSS IN1 dantenna A=35.0028 P=58.08 m=2
* device instance $3063 r0 *1 1195.06,1000 dantenna
D$3063 VSS OUT1 dantenna A=35.0028 P=58.08 m=2
* device instance $3065 r0 *1 222.54,1017.63 dantenna
D$3065 VSS \$1969 dantenna A=1.984 P=7.48 m=1
* device instance $3066 r0 *1 417.63,1077.46 dantenna
D$3066 VSS \$1718 dantenna A=1.984 P=7.48 m=1
* device instance $3067 r0 *1 517.63,1077.46 dantenna
D$3067 VSS \$2028 dantenna A=1.984 P=7.48 m=1
* device instance $3068 r0 *1 705.225,1077.46 dantenna
D$3068 VSS \$2013 dantenna A=1.984 P=7.48 m=1
* device instance $3069 r0 *1 805.225,1077.46 dantenna
D$3069 VSS \$2014 dantenna A=1.984 P=7.48 m=1
* device instance $3070 r0 *1 905.225,1077.46 dantenna
D$3070 VSS \$2015 dantenna A=1.984 P=7.48 m=1
* device instance $3071 r0 *1 664.54,1195.81 dantenna
D$3071 VSS CK3 dantenna A=35.0028 P=58.08 m=2
* device instance $3073 r0 *1 764.54,1195.81 dantenna
D$3073 VSS CK2 dantenna A=35.0028 P=58.08 m=2
* device instance $3075 r0 *1 864.54,1195.81 dantenna
D$3075 VSS CK1 dantenna A=35.0028 P=58.08 m=2
* device instance $3077 r0 *1 264.765,1192.65 dantenna
D$3077 VSS \$2089 dantenna A=0.192 P=1.88 m=1
* device instance $3078 r0 *1 400,1195.06 dantenna
D$3078 VSS VREF dantenna A=35.0028 P=58.08 m=2
* device instance $3079 r0 *1 500,1195.06 dantenna
D$3079 VSS VLDO dantenna A=35.0028 P=58.08 m=2
* device instance $3080 r0 *1 564.765,1192.65 dantenna
D$3080 VSS \$2090 dantenna A=0.192 P=1.88 m=1
* device instance $3081 r0 *1 964.765,1192.65 dantenna
D$3081 VSS \$2091 dantenna A=0.192 P=1.88 m=1
* device instance $3084 r0 *1 264.54,163.19 dpantenna
D$3084 VSS AVDD dpantenna A=35.0028 P=58.08 m=4
* device instance $3088 r0 *1 464.54,163.19 dpantenna
D$3088 RES IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3090 r0 *1 564.54,163.19 dpantenna
D$3090 VSS IOVDD dpantenna A=35.0028 P=58.08 m=6
* device instance $3092 r0 *1 664.54,163.19 dpantenna
D$3092 CK4 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3094 r0 *1 764.54,163.19 dpantenna
D$3094 CK5 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3096 r0 *1 864.54,163.19 dpantenna
D$3096 CK6 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3100 r0 *1 227.51,315.46 dpantenna
D$3100 \$288 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3101 r0 *1 227.51,415.46 dpantenna
D$3101 \$403 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3102 r0 *1 227.51,515.46 dpantenna
D$3102 \$587 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3103 r0 *1 227.51,615.46 dpantenna
D$3103 \$953 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3104 r0 *1 227.51,715.46 dpantenna
D$3104 \$1218 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3105 r0 *1 227.51,815.46 dpantenna
D$3105 \$1344 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3106 r0 *1 227.51,915.46 dpantenna
D$3106 \$1854 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3107 r0 *1 227.51,1015.46 dpantenna
D$3107 \$1969 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3108 r0 *1 415.46,1072.49 dpantenna
D$3108 \$1718 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3109 r0 *1 515.46,1072.49 dpantenna
D$3109 \$2028 AVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3110 r0 *1 503.055,227.51 dpantenna
D$3110 \$129 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3111 r0 *1 703.055,227.51 dpantenna
D$3111 \$130 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3112 r0 *1 803.055,227.51 dpantenna
D$3112 \$132 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3113 r0 *1 903.055,227.51 dpantenna
D$3113 \$133 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3114 r0 *1 703.055,1072.49 dpantenna
D$3114 \$2013 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3115 r0 *1 803.055,1072.49 dpantenna
D$3115 \$2014 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3116 r0 *1 903.055,1072.49 dpantenna
D$3116 \$2015 IOVDD dpantenna A=3.1872 P=11.24 m=1
* device instance $3117 r0 *1 1138.81,277.975 dpantenna
D$3117 \$216 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $3118 r0 *1 135.96,300 dpantenna
D$3118 IN6 AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3120 r0 *1 1159.54,300 dpantenna
D$3120 OUT6 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3122 r0 *1 135.96,400 dpantenna
D$3122 IN5 AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3124 r0 *1 1138.81,377.975 dpantenna
D$3124 \$331 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $3125 r0 *1 1159.54,400 dpantenna
D$3125 OUT5 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3127 r0 *1 135.96,500 dpantenna
D$3127 IN4 AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3129 r0 *1 1138.81,477.975 dpantenna
D$3129 \$446 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $3130 r0 *1 1159.54,500 dpantenna
D$3130 OUT4 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3132 r0 *1 135.96,600 dpantenna
D$3132 VLO AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3136 r0 *1 135.96,700 dpantenna
D$3136 VHI AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3138 r0 *1 1138.81,777.975 dpantenna
D$3138 \$1272 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $3139 r0 *1 135.96,800 dpantenna
D$3139 IN3 AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3141 r0 *1 1159.54,800 dpantenna
D$3141 OUT3 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3143 r0 *1 135.96,900 dpantenna
D$3143 IN2 AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3145 r0 *1 1138.81,877.975 dpantenna
D$3145 \$1712 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $3146 r0 *1 1159.54,900 dpantenna
D$3146 OUT2 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3148 r0 *1 135.96,1000 dpantenna
D$3148 IN1 AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3150 r0 *1 1138.81,977.975 dpantenna
D$3150 \$1897 IOVDD dpantenna A=0.192 P=1.88 m=1
* device instance $3151 r0 *1 1159.54,1000 dpantenna
D$3151 OUT1 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3153 r0 *1 664.54,1136.81 dpantenna
D$3153 CK3 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3155 r0 *1 764.54,1136.81 dpantenna
D$3155 CK2 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3157 r0 *1 864.54,1136.81 dpantenna
D$3157 CK1 IOVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3159 r0 *1 400,1159.54 dpantenna
D$3159 VREF AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3161 r0 *1 500,1159.54 dpantenna
D$3161 VLDO AVDD dpantenna A=35.0028 P=58.08 m=2
* device instance $3163 r0 *1 500.685,221.11 rppd
R$3163 RES \$129 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3164 r0 *1 700.685,221.11 rppd
R$3164 CK4 \$130 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3165 r0 *1 800.685,221.11 rppd
R$3165 CK5 \$132 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3166 r0 *1 900.685,221.11 rppd
R$3166 CK6 \$133 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3167 r0 *1 88.75,326.305 rppd
R$3167 VSS \$225 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $3168 r0 *1 147.75,326.305 rppd
R$3168 AVDD \$226 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $3169 r0 *1 221.11,313.09 rppd
R$3169 IN6 \$288 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3170 r0 *1 88.75,426.305 rppd
R$3170 VSS \$340 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $3171 r0 *1 147.75,426.305 rppd
R$3171 AVDD \$341 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $3172 r0 *1 221.11,413.09 rppd
R$3172 IN5 \$403 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3173 r0 *1 88.75,526.305 rppd
R$3173 VSS \$455 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $3174 r0 *1 147.75,526.305 rppd
R$3174 AVDD \$456 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $3175 r0 *1 221.11,513.09 rppd
R$3175 IN4 \$587 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3176 r0 *1 88.75,626.305 rppd
R$3176 VSS \$845 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $3177 r0 *1 147.75,626.305 rppd
R$3177 AVDD \$846 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $3178 r0 *1 221.11,613.09 rppd
R$3178 VLO \$953 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3179 r0 *1 1161.29,678.875 rppd
R$3179 IOVDD \$1185 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $3180 r0 *1 221.11,713.09 rppd
R$3180 VHI \$1218 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3181 r0 *1 88.75,726.305 rppd
R$3181 VSS \$1190 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $3182 r0 *1 147.75,726.305 rppd
R$3182 AVDD \$1191 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $3183 r0 *1 88.75,826.305 rppd
R$3183 VSS \$1282 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $3184 r0 *1 147.75,826.305 rppd
R$3184 AVDD \$1283 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $3185 r0 *1 221.11,813.09 rppd
R$3185 IN3 \$1344 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3186 r0 *1 221.11,913.09 rppd
R$3186 IN2 \$1854 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3187 r0 *1 88.75,926.305 rppd
R$3187 VSS \$1736 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $3188 r0 *1 147.75,926.305 rppd
R$3188 AVDD \$1737 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $3189 r0 *1 88.75,1026.305 rppd
R$3189 VSS \$1906 rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $3190 r0 *1 147.75,1026.305 rppd
R$3190 AVDD \$1907 rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $3191 r0 *1 221.11,1013.09 rppd
R$3191 IN1 \$1969 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3192 r0 *1 413.09,1076.03 rppd
R$3192 \$1718 VREF rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3193 r0 *1 513.09,1076.03 rppd
R$3193 \$2028 VLDO rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3194 r0 *1 700.685,1076.03 rppd
R$3194 \$2013 CK3 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3195 r0 *1 800.685,1076.03 rppd
R$3195 \$2014 CK2 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3196 r0 *1 900.685,1076.03 rppd
R$3196 \$2015 CK1 rppd w=1 l=2 ps=0 b=0 m=1
* device instance $3197 r0 *1 278.875,1161.29 rppd
R$3197 AVDD \$2148 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $3198 r0 *1 426.305,1138.49 rppd
R$3198 \$2106 AVDD rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $3199 r0 *1 526.305,1138.49 rppd
R$3199 \$2107 AVDD rppd w=0.5 l=12.9 ps=0 b=0 m=1
* device instance $3200 r0 *1 578.875,1161.29 rppd
R$3200 IOVDD \$2149 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $3201 r0 *1 978.875,1161.29 rppd
R$3201 VDD \$2150 rppd w=1 l=0 ps=0 b=25 m=1
* device instance $3202 r0 *1 426.305,1206.85 rppd
R$3202 \$2220 VSS rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $3203 r0 *1 526.305,1206.85 rppd
R$3203 \$2221 VSS rppd w=0.5 l=3.54 ps=0 b=0 m=1
* device instance $3204 r0 *1 506.575,859.565 rhigh
R$3204 VSS \$1621 rhigh w=0.5 l=0.96 ps=0 b=0 m=2
* device instance $3208 r0 *1 543.535,883.575 rhigh
R$3208 \$1377 \$1378 rhigh w=0.5 l=3.84 ps=0 b=0 m=1
* device instance $3210 r0 *1 430.19,624.19 cap_cmim
C$3210 \$1071 \$1016 cap_cmim w=8.16 l=8.16 m=1
* device instance $3211 r0 *1 479.935,615.55 cap_cmim
C$3211 \$994 \$1017 cap_cmim w=5.77 l=5.77 m=1
* device instance $3212 r0 *1 443.88,615.55 cap_cmim
C$3212 \$993 \$1015 cap_cmim w=5.77 l=5.77 m=1
* device instance $3213 r0 *1 509.38,615.465 cap_cmim
C$3213 \$1061 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $3214 r0 *1 485.88,542.236 cap_cmim
C$3214 \$564 \$798 cap_cmim w=8.16 l=8.16 m=1
* device instance $3215 r0 *1 439.56,542.231 cap_cmim
C$3215 \$757 \$789 cap_cmim w=8.16 l=8.16 m=1
* device instance $3216 r0 *1 597.775,848.635 cap_cmim
C$3216 \$1421 \$1418 cap_cmim w=5.77 l=5.77 m=1
* device instance $3217 r0 *1 576.185,848.635 cap_cmim
C$3217 \$1420 \$1417 cap_cmim w=5.77 l=5.77 m=1
* device instance $3218 r0 *1 430.955,540.411 cap_cmim
C$3218 \$789 \$791 cap_cmim w=5.77 l=5.77 m=1
* device instance $3219 r0 *1 597.895,835.415 cap_cmim
C$3219 \$1387 \$1421 cap_cmim w=8.16 l=8.16 m=1
* device instance $3220 r0 *1 466.245,624.19 cap_cmim
C$3220 \$1072 \$1018 cap_cmim w=8.16 l=8.16 m=1
* device instance $3221 r0 *1 477.165,625.165 cap_cmim
C$3221 \$1106 \$994 cap_cmim w=8.16 l=8.16 m=1
* device instance $3222 r0 *1 576.305,835.415 cap_cmim
C$3222 \$1386 \$1420 cap_cmim w=8.16 l=8.16 m=1
* device instance $3223 r0 *1 441.11,625.165 cap_cmim
C$3223 \$1105 \$993 cap_cmim w=8.16 l=8.16 m=1
* device instance $3224 r0 *1 609.13,835.275 cap_cmim
C$3224 \$1383 \$1391 cap_cmim w=8.16 l=8.16 m=1
* device instance $3225 r0 *1 587.54,835.275 cap_cmim
C$3225 \$1382 \$1406 cap_cmim w=8.16 l=8.16 m=1
* device instance $3226 r0 *1 623.755,834.77 cap_cmim
C$3226 \$1384 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $3227 r0 *1 450.88,542.236 cap_cmim
C$3227 \$752 \$797 cap_cmim w=8.16 l=8.16 m=1
* device instance $3228 r0 *1 474.56,542.231 cap_cmim
C$3228 \$758 \$790 cap_cmim w=8.16 l=8.16 m=1
* device instance $3229 r0 *1 429.41,682.847 cap_cmim
C$3229 VSS VLDO cap_cmim w=140 l=225 m=1
* device instance $3230 r0 *1 429.41,826.865 cap_cmim
C$3230 \$1378 VLDO cap_cmim w=60 l=60 m=1
* device instance $3231 r0 *1 473.164,512.175 cap_cmim
C$3231 \$565 VSS cap_cmim w=5.77 l=5.77 m=1
* device instance $3232 r0 *1 465.955,540.411 cap_cmim
C$3232 \$790 \$792 cap_cmim w=5.77 l=5.77 m=1
.ENDS UHEE628_S2024

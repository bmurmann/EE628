** sch_path: /foss/designs/comp_5_split2.sch
.subckt comp_5_split2 VDD out1p out2m out1m VSS
*.PININFO out1m:B out2m:B out1p:B VSS:B VDD:B
M3 out2m out1m VDD VDD sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M12 out2m out1p VDD VDD sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M15 out2m out1p net1 VSS sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M16 net1 out1m VSS VSS sg13_lv_nmos L=0.13u W=2u ng=1 m=1
.ends
.end

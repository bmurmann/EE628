* Extracted by KLayout with SG13G2 LVS runset on : 01/05/2024 21:50

* cell sg13g2_IOPadInOut16mA
.SUBCKT sg13g2_IOPadInOut16mA
* net 5 sub!
* net 7 dant
* net 10 PAD
* net 11 sub!
* net 12 dant
* net 14 diodevss_4kv
* net 15 dant
* net 20 sub!
* net 21 PAD
* net 24 dpant
* net 25 diodevdd_4kv
* net 26 dpant
* net 30 sub!
* net 33 dpant
* net 39 PAD
* net 40 sub!
* net 41 rppd r=793.834
* net 42 IOVSS
* net 43 sub!
* net 45 dant
* net 46 IOVDD
* net 48 dpant
* net 50 CORE
* net 102 sub!
* device instance $1 r0 *1 18.685,171.175 sg13_lv_nmos
M$1 102 87 58 102 sg13_lv_nmos W=3.9299999999999993 L=0.12999999999999998
* device instance $2 r0 *1 19.195,171.175 sg13_lv_nmos
M$2 58 88 102 102 sg13_lv_nmos W=3.9299999999999993 L=0.12999999999999998
* device instance $3 r0 *1 60.255,159.005 sg13_lv_nmos
M$3 67 69 102 102 sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $4 r0 *1 23.485,171.175 sg13_lv_nmos
M$4 102 89 88 102 sg13_lv_nmos W=3.9299999999999993 L=0.12999999999999998
* device instance $5 r0 *1 18.685,159.005 sg13_lv_nmos
M$5 57 58 102 102 sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $6 r0 *1 22.195,159.005 sg13_lv_nmos
M$6 59 60 102 102 sg13_lv_nmos W=2.7499999999999996 L=0.12999999999999995
* device instance $7 r0 *1 21.085,171.175 sg13_lv_nmos
M$7 102 87 91 102 sg13_lv_nmos W=3.9299999999999993 L=0.12999999999999998
* device instance $8 r0 *1 21.595,171.175 sg13_lv_nmos
M$8 91 89 60 102 sg13_lv_nmos W=3.9299999999999993 L=0.12999999999999998
* device instance $9 r0 *1 61.765,159.055 sg13_hv_nmos
M$9 102 38 69 102 sg13_hv_nmos W=2.6499999999999995 L=0.4499999999999999
* device instance $10 r0 *1 18.845,155.32 sg13_hv_nmos
M$10 51 57 102 102 sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $11 r0 *1 19.675,155.32 sg13_hv_nmos
M$11 102 58 52 102 sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $12 r0 *1 34.58,10.95 sg13_hv_nmos
M$12 102 6 1 102 sg13_hv_nmos W=35.199999999999996 L=0.5999999999999998
* device instance $20 r0 *1 24.525,155.32 sg13_hv_nmos
M$20 102 54 32 102 sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $21 r0 *1 21.015,155.32 sg13_hv_nmos
M$21 102 52 6 102 sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $22 r0 *1 22.355,155.32 sg13_hv_nmos
M$22 53 59 102 102 sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $23 r0 *1 23.185,155.32 sg13_hv_nmos
M$23 102 60 54 102 sg13_hv_nmos W=1.8999999999999997 L=0.4499999999999999
* device instance $24 r0 *1 18.685,176.585 sg13_lv_pmos
M$24 37 87 97 37 sg13_lv_pmos W=4.409999999999999 L=0.12999999999999995
* device instance $25 r0 *1 19.195,176.585 sg13_lv_pmos
M$25 97 88 58 37 sg13_lv_pmos W=4.409999999999999 L=0.12999999999999995
* device instance $26 r0 *1 22.195,163.995 sg13_lv_pmos
M$26 59 60 37 37 sg13_lv_pmos W=4.749999999999999 L=0.12999999999999998
* device instance $27 r0 *1 21.085,176.585 sg13_lv_pmos
M$27 37 87 60 37 sg13_lv_pmos W=4.409999999999999 L=0.12999999999999995
* device instance $28 r0 *1 21.595,176.585 sg13_lv_pmos
M$28 60 89 37 37 sg13_lv_pmos W=4.409999999999999 L=0.12999999999999995
* device instance $29 r0 *1 18.685,163.995 sg13_lv_pmos
M$29 57 58 37 37 sg13_lv_pmos W=4.749999999999999 L=0.12999999999999998
* device instance $30 r0 *1 60.255,163.995 sg13_lv_pmos
M$30 67 69 37 37 sg13_lv_pmos W=4.749999999999999 L=0.12999999999999998
* device instance $31 r0 *1 23.485,176.585 sg13_lv_pmos
M$31 37 89 88 37 sg13_lv_pmos W=4.409999999999999 L=0.12999999999999995
* device instance $32 r0 *1 61.765,163.945 sg13_hv_pmos
M$32 37 38 69 37 sg13_hv_pmos W=4.6499999999999995 L=0.44999999999999984
* device instance $33 r0 *1 24.525,151.18 sg13_hv_pmos
M$33 36 54 32 36 sg13_hv_pmos W=3.899999999999999 L=0.4499999999999999
* device instance $34 r0 *1 21.015,151.18 sg13_hv_pmos
M$34 36 52 6 36 sg13_hv_pmos W=3.899999999999999 L=0.4499999999999999
* device instance $35 r0 *1 22.355,151.18 sg13_hv_pmos
M$35 53 54 36 36 sg13_hv_pmos W=0.29999999999999993 L=0.44999999999999984
* device instance $36 r0 *1 23.185,151.18 sg13_hv_pmos
M$36 36 53 54 36 sg13_hv_pmos W=0.29999999999999993 L=0.44999999999999984
* device instance $37 r0 *1 18.845,151.18 sg13_hv_pmos
M$37 51 52 36 36 sg13_hv_pmos W=0.29999999999999993 L=0.44999999999999984
* device instance $38 r0 *1 19.675,151.18 sg13_hv_pmos
M$38 36 51 52 36 sg13_hv_pmos W=0.29999999999999993 L=0.44999999999999984
* device instance $39 r0 *1 34.58,78.18 sg13_hv_pmos
M$39 22 32 1 22 sg13_hv_pmos W=106.55999999999996 L=0.5999999999999999
* device instance $55 r0 *1 17.975,12.83 dantenna
D$55 102 6 dantenna A=0.192 P=1.88 m=1
* device instance $56 r0 *1 40,20.44 dantenna
D$56 102 1 dantenna A=35.0028 P=58.08 m=2
* device instance $58 r0 *1 65.225,142.54 dantenna
D$58 102 38 dantenna A=1.984 P=7.48 m=1
* device instance $59 r0 *1 40,55.96 dpantenna
D$59 1 22 dpantenna A=35.0028 P=58.08 m=2
* device instance $61 r0 *1 17.975,81.19 dpantenna
D$61 32 22 dpantenna A=0.192 P=1.88 m=1
* device instance $62 r0 *1 63.055,147.51 dpantenna
D$62 38 36 dpantenna A=3.1872 P=11.24 m=1
* device instance $63 r0 *1 60.685,141.11 res_rppd
R$63 1 38 res_rppd w=0.9999999999999998 l=1.9999999999999996 b=0.0 ps=0.0 m=1.0
.ENDS sg13g2_IOPadInOut16mA

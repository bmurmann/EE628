* Extracted by KLayout with SG13G2 LVS runset on : 09/05/2024 08:44

* cell comp_5_splitTop1
* pin sub!
.SUBCKT comp_5_splitTop1 sub!
* device instance $1 r0 *1 -6.53,-4.181 sg13_lv_nmos
M$1 sub! \$8 \$2 sub! sg13_lv_nmos W=2.0 L=1.0
* device instance $2 r0 *1 -3.17,-2.514 sg13_lv_nmos
M$2 \$4 \$23 \$9 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $3 r0 *1 -1.525,-2.514 sg13_lv_nmos
M$3 \$9 \$16 \$2 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $4 r0 *1 -6.53,1.48 sg13_lv_nmos
M$4 sub! \$27 \$15 sub! sg13_lv_nmos W=2.0 L=1.0
* device instance $5 r0 *1 -3.17,3.147 sg13_lv_nmos
M$5 \$23 \$4 \$28 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $6 r0 *1 -1.525,3.147 sg13_lv_nmos
M$6 \$28 \$16 \$15 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $7 r0 *1 -5.021,-3.488 sg13_lv_pmos
M$7 \$3 \$23 \$4 \$3 sg13_lv_pmos W=4.0 L=0.13
* device instance $8 r0 *1 0.326,-3.488 sg13_lv_pmos
M$8 \$4 \$16 \$3 \$3 sg13_lv_pmos W=4.0 L=0.13
* device instance $9 r0 *1 -5.021,2.173 sg13_lv_pmos
M$9 \$3 \$4 \$23 \$3 sg13_lv_pmos W=4.0 L=0.13
* device instance $10 r0 *1 0.326,2.173 sg13_lv_pmos
M$10 \$23 \$16 \$3 \$3 sg13_lv_pmos W=4.0 L=0.13
.ENDS comp_5_splitTop1

* Extracted by KLayout with SG13G2 LVS runset on : 09/05/2024 15:26

* cell Team5_split1
* pin sub!
.SUBCKT Team5_split1 sub!
* device instance $1 r0 *1 -15.942,-16.032 sg13_lv_nmos
M$1 \$7 \$8 sub! sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $2 r0 *1 -15.432,-15.982 sg13_lv_nmos
M$2 sub! \$9 \$17 sub! sg13_lv_nmos W=0.64 L=0.13
* device instance $3 r0 *1 -14.922,-15.982 sg13_lv_nmos
M$3 \$17 \$47 \$8 sub! sg13_lv_nmos W=0.64 L=0.13
* device instance $4 r0 *1 -3.802,-15.982 sg13_lv_nmos
M$4 \$11 \$10 \$16 sub! sg13_lv_nmos W=0.64 L=0.13
* device instance $5 r0 *1 -3.292,-15.982 sg13_lv_nmos
M$5 sub! \$12 \$16 sub! sg13_lv_nmos W=0.64 L=0.13
* device instance $6 r0 *1 -2.782,-16.032 sg13_lv_nmos
M$6 sub! \$11 \$13 sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $7 r0 *1 -20.688,-15.088 sg13_lv_nmos
M$7 \$3 \$7 \$20 sub! sg13_lv_nmos W=0.5 L=0.13
* device instance $8 r0 *1 1.964,-15.088 sg13_lv_nmos
M$8 \$3 \$13 \$38 sub! sg13_lv_nmos W=0.5 L=0.13
* device instance $9 r0 *1 -21.845,-10.363 sg13_lv_nmos
M$9 \$20 \$10 \$37 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $10 r0 *1 3.121,-10.363 sg13_lv_nmos
M$10 \$110 \$47 \$38 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $11 r0 *1 -36.647,-6.47 sg13_lv_nmos
M$11 \$91 \$47 \$1 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $12 r0 *1 -32.071,-6.47 sg13_lv_nmos
M$12 \$1 \$48 \$50 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $13 r0 *1 13.347,-6.47 sg13_lv_nmos
M$13 \$51 \$49 \$5 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $14 r0 *1 17.923,-6.47 sg13_lv_nmos
M$14 \$5 \$10 \$92 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $15 r0 *1 -21.45,-3.88 sg13_lv_nmos
M$15 sub! \$10 \$28 sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $16 r0 *1 -18.102,-3.785 sg13_lv_nmos
M$16 sub! \$9 \$64 sub! sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $17 r0 *1 -17.252,-3.88 sg13_lv_nmos
M$17 sub! \$47 \$72 sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $18 r0 *1 -16.942,-3.88 sg13_lv_nmos
M$18 \$72 \$64 \$65 sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $19 r0 *1 -1.782,-3.88 sg13_lv_nmos
M$19 \$67 \$68 \$73 sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $20 r0 *1 -1.472,-3.88 sg13_lv_nmos
M$20 \$73 \$10 sub! sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $21 r0 *1 -0.622,-3.785 sg13_lv_nmos
M$21 sub! \$12 \$68 sub! sg13_lv_nmos W=0.55 L=0.12999999999999998
* device instance $22 r0 *1 2.726,-3.88 sg13_lv_nmos
M$22 \$30 \$47 sub! sub! sg13_lv_nmos W=0.74 L=0.13
* device instance $23 r0 *1 -26.132,1.508 sg13_lv_nmos
M$23 \$50 \$50 sub! sub! sg13_lv_nmos W=2.5 L=1.5
* device instance $24 r0 *1 7.408,1.508 sg13_lv_nmos
M$24 sub! \$51 \$51 sub! sg13_lv_nmos W=2.5 L=1.5
* device instance $25 r0 *1 -26.132,11.054 sg13_lv_nmos
M$25 \$110 \$4 sub! sub! sg13_lv_nmos W=2.5 L=1.5
* device instance $26 r0 *1 7.408,11.054 sg13_lv_nmos
M$26 sub! \$6 \$109 sub! sg13_lv_nmos W=2.5 L=1.5
* device instance $27 r0 *1 -21.194,13.511 sg13_lv_nmos
M$27 \$110 \$113 \$91 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $28 r0 *1 -16.618,13.511 sg13_lv_nmos
M$28 \$91 \$10 \$4 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $29 r0 *1 -2.106,13.511 sg13_lv_nmos
M$29 \$6 \$47 \$92 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $30 r0 *1 2.47,13.511 sg13_lv_nmos
M$30 \$92 \$113 \$109 sub! sg13_lv_nmos W=2.0 L=0.13
* device instance $31 r0 *1 -15.942,-14.482 sg13_lv_pmos
M$31 \$7 \$8 \$21 \$21 sg13_lv_pmos W=1.12 L=0.13
* device instance $32 r0 *1 -15.432,-14.342 sg13_lv_pmos
M$32 \$21 \$9 \$8 \$21 sg13_lv_pmos W=0.84 L=0.13
* device instance $33 r0 *1 -14.922,-14.342 sg13_lv_pmos
M$33 \$8 \$47 \$21 \$21 sg13_lv_pmos W=0.84 L=0.13
* device instance $34 r0 *1 -3.802,-14.342 sg13_lv_pmos
M$34 \$21 \$10 \$11 \$21 sg13_lv_pmos W=0.84 L=0.13
* device instance $35 r0 *1 -3.292,-14.342 sg13_lv_pmos
M$35 \$21 \$12 \$11 \$21 sg13_lv_pmos W=0.84 L=0.13
* device instance $36 r0 *1 -2.782,-14.482 sg13_lv_pmos
M$36 \$21 \$11 \$13 \$21 sg13_lv_pmos W=1.12 L=0.13
* device instance $37 r0 *1 -16.213,-10.361 sg13_lv_pmos
M$37 \$20 \$28 \$37 \$29 sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $41 r0 *1 -4.041,-10.361 sg13_lv_pmos
M$41 \$38 \$30 \$110 \$29 sg13_lv_pmos W=6.0 L=0.12999999999999998
* device instance $45 r0 *1 -13.991,-2.732 sg13_lv_pmos
M$45 \$66 \$65 \$20 \$29 sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $46 r0 *1 -4.733,-2.732 sg13_lv_pmos
M$46 \$38 \$67 \$66 \$29 sg13_lv_pmos W=1.5 L=0.12999999999999998
* device instance $47 r0 *1 -18.102,-2.36 sg13_lv_pmos
M$47 \$64 \$9 \$21 \$21 sg13_lv_pmos W=0.84 L=0.13
* device instance $48 r0 *1 -17.562,-2.22 sg13_lv_pmos
M$48 \$21 \$47 \$65 \$21 sg13_lv_pmos W=1.12 L=0.13
* device instance $49 r0 *1 -17.052,-2.22 sg13_lv_pmos
M$49 \$65 \$64 \$21 \$21 sg13_lv_pmos W=1.12 L=0.13
* device instance $50 r0 *1 -0.622,-2.36 sg13_lv_pmos
M$50 \$21 \$12 \$68 \$21 sg13_lv_pmos W=0.84 L=0.13
* device instance $51 r0 *1 -1.672,-2.22 sg13_lv_pmos
M$51 \$21 \$68 \$67 \$21 sg13_lv_pmos W=1.12 L=0.13
* device instance $52 r0 *1 -1.162,-2.22 sg13_lv_pmos
M$52 \$67 \$10 \$21 \$21 sg13_lv_pmos W=1.12 L=0.13
* device instance $53 r0 *1 -21.44,-2.205 sg13_lv_pmos
M$53 \$21 \$10 \$28 \$21 sg13_lv_pmos W=1.12 L=0.13
* device instance $54 r0 *1 2.716,-2.205 sg13_lv_pmos
M$54 \$30 \$47 \$21 \$21 sg13_lv_pmos W=1.12 L=0.13
* device instance $55 r0 *1 -38.19,1.524 sg13_lv_pmos
M$55 \$50 \$50 \$29 \$29 sg13_lv_pmos W=10.0 L=1.5
* device instance $59 r0 *1 13.826,1.524 sg13_lv_pmos
M$59 \$51 \$51 \$29 \$29 sg13_lv_pmos W=10.0 L=1.5
* device instance $63 r0 *1 -38.19,11.07 sg13_lv_pmos
M$63 \$110 \$4 \$29 \$29 sg13_lv_pmos W=10.0 L=1.5
* device instance $67 r0 *1 13.826,11.07 sg13_lv_pmos
M$67 \$109 \$6 \$29 \$29 sg13_lv_pmos W=10.0 L=1.5
* device instance $71 r0 *1 5.01,-18.47 cap_cmim
C$71 \$5 \$38 cap_cmim w=5.77 l=5.77 m=1
* device instance $72 r0 *1 -40.279,-18.475 cap_cmim
C$72 \$4 \$1 cap_cmim w=8.16 l=8.16 m=1
* device instance $73 r0 *1 -30.704,-18.47 cap_cmim
C$73 \$1 \$20 cap_cmim w=5.77 l=5.77 m=1
* device instance $74 r0 *1 12.195,-18.475 cap_cmim
C$74 \$6 \$5 cap_cmim w=8.16 l=8.16 m=1
* device instance $75 r0 *1 -22.46,1.213 cap_cmim
C$75 \$91 \$110 cap_cmim w=8.16 l=8.16 m=1
* device instance $76 r0 *1 -5.624,1.213 cap_cmim
C$76 \$92 \$109 cap_cmim w=8.16 l=8.16 m=1
.ENDS Team5_split1

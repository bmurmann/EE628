** sch_path: /foss/designs/EE628/5_Design/3_Real_circuits/tb_UHEE628_S2024.sch
**.subckt tb_UHEE628_S2024
x1 net1 ck1 ck3 vdd ck2 vdd GND out1 GND GND out2 out3 GND iovdd vhi vlo out4 GND out5 GND out6 GND ck6 ck5 ck4 reset GND
+ UHEE628_S2024
V1 iovdd GND 3
V2 vdd GND 1.2
* noconn #net1
V3 vlo GND 0.3
V4 vhi GND 0.9
C1 out6 GND 1p m=1
C2 out5 GND 1p m=1
C3 out4 GND 1p m=1
C4 out3 GND 1p m=1
C5 out2 GND 1p m=1
C6 out1 GND 1p m=1
* noconn ck1
* noconn ck3
* noconn ck2
* noconn ck6
* noconn ck5
* noconn ck4
* noconn reset
**** begin user architecture code



* ngspice commands
.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt
.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ
.inc /foss/pdks/sg13g2/libs.tech/ngspice/models/diodes.lib
.inc "../../4_Layout/Team 1/Team1_sim.spice"
.inc "../../4_Layout/Team 2 - Transformer Monster Tractors/Team_2_sim.spice"
.inc "../../4_Layout/Team 3/Team3_sim.spice"
.inc "../../4_Layout/Team 4/Team4_sim.spice"
.inc "../../4_Layout/Team 5/Team5_sim.spice"
.inc "../../4_Layout/Team 6/Team6_sim.spice"
.inc "../stimulus_gen/inc_clocks.spice"
.inc ../sg13g2_stdcell.spice
.inc ../sg13g2_io.spi
.options gmin=1e-8 keepopinfo

.control
optran 0 0 0 100p 2n 0
op
tran 1u 250u
plot reset ck1
plot out1 out2
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/EE628/5_Design/3_Real_circuits/UHEE628_S2024.sym # of pins=27
** sym_path: /foss/designs/EE628/5_Design/3_Real_circuits/UHEE628_S2024.sym
** sch_path: /foss/designs/EE628/5_Design/3_Real_circuits/UHEE628_S2024.sch
.subckt UHEE628_S2024 vldo ck1 ck3 avdd ck2 VDD vref out1 in1 in2 out2 out3 in3 iovdd vhi vlo out4 in4 out5 in5 out6 in6 ck6 ck5
+ ck4 res VSS
*.ipin in1
*.ipin in2
*.ipin in3
*.ipin in4
*.ipin in5
*.ipin in6
*.iopin iovdd
*.iopin vlo
*.iopin avdd
*.opin out1
*.opin out2
*.opin out3
*.opin out4
*.opin out5
*.opin out6
*.iopin VSS
*.iopin VDD
*.iopin vldo
*.ipin ck3
*.ipin ck2
*.ipin ck1
*.ipin vref
*.ipin res
*.ipin ck4
*.ipin ck5
*.ipin ck6
*.iopin vhi
x10 vref ck3 vldo ck1 ck2 ck1_c ck3_c vref_c ck2_c out1_c in1 out1 in2 out2 out2_c in2_c VDD out3 in3_c in3 out3_c avdd iovdd vhi
+ vlo out4 in4_c in4 out4_c out5 in5_c out5_c in5 in6 in6_c out6 out6_c ck5_c ck4_c res_c ck6_c ck6 ck5 ck4 res in1_c VSS padring
x1 vhi vlo avdd VSS in1_c out1_c res_c ck1_c Team1
x2 vlo vhi vldo VSS iovdd vref_c in2_c out2_c res_c ck2_c Team_2
x4 vhi vlo avdd VSS in4_c out4_c res_c ck4_c Team4
x5 vhi vlo avdd VSS in5_c out5_c res_c ck5_c Team5
x6 vhi vlo avdd VSS in6_c out6_c res_c ck6_c Team6
x7 vhi vlo avdd VSS in3_c out3_c res_c ck3_c Team3
.ends


* expanding   symbol:  padring.sym # of pins=47
** sym_path: /foss/designs/EE628/5_Design/3_Real_circuits/padring.sym
** sch_path: /foss/designs/EE628/5_Design/3_Real_circuits/padring.sch
.subckt padring vref ck3 vldo ck1 ck2 ck1_c ck3_c vref_c ck2_c out1_c in1 out1 in2 out2 out2_c in2_c vdd out3 in3_c in3 out3_c
+ avdd iovdd vhi vlo out4 in4_c in4 out4_c out5 in5_c out5_c in5 in6 in6_c out6 out6_c ck5_c ck4_c res_c ck6_c ck6 ck5 ck4 res in1_c vss
*.ipin in1
*.ipin in2
*.ipin in3
*.iopin vhi
*.iopin vlo
*.ipin in4
*.ipin in5
*.ipin in6
*.opin out1
*.opin out2
*.opin out3
*.opin out4
*.opin out5
*.opin out6
*.ipin res
*.ipin ck4
*.ipin ck5
*.ipin ck6
*.ipin vref
*.ipin ck3
*.ipin ck2
*.ipin ck1
*.opin in1_c
*.opin in2_c
*.opin in3_c
*.opin in4_c
*.opin in5_c
*.opin in6_c
*.opin res_c
*.opin ck4_c
*.opin ck5_c
*.opin ck6_c
*.ipin out1_c
*.ipin out2_c
*.ipin out3_c
*.ipin out4_c
*.ipin out5_c
*.ipin out6_c
*.opin vref_c
*.opin ck3_c
*.opin ck2_c
*.opin ck1_c
*.iopin vldo
*.iopin avdd
*.iopin vss
*.iopin iovdd
*.iopin vdd
xp1 vss avdd vss avdd in1 in1_c sg13g2_IOPadAnalog
xp26 vss vdd vss iovdd ck1_c ck1 sg13g2_IOPadIn
xp24 vss vdd vss iovdd out1_c out1 sg13g2_IOPadOut16mA
xp32 vss avdd vss avdd sg13g2_IOPadVdd
xp9 vss avdd vss avdd sg13g2_IOPadVss
xp2 vss avdd vss avdd in2 in2_c sg13g2_IOPadAnalog
xp3 vss avdd vss avdd in3 in3_c sg13g2_IOPadAnalog
xp4 vss avdd vss avdd vhi net1 sg13g2_IOPadAnalog
xp5 vss avdd vss avdd vlo net2 sg13g2_IOPadAnalog
xp6 vss avdd vss avdd in4 in4_c sg13g2_IOPadAnalog
xp7 vss avdd vss avdd in5 in5_c sg13g2_IOPadAnalog
xp8 vss avdd vss avdd in6 in6_c sg13g2_IOPadAnalog
xp23 vss vdd vss iovdd out2_c out2 sg13g2_IOPadOut16mA
xp22 vss vdd vss iovdd out3_c out3 sg13g2_IOPadOut16mA
xp21 vss vdd vss iovdd sg13g2_IOPadIOVdd
xp20 vss vdd vss iovdd sg13g2_IOPadIOVss
xp19 vss vdd vss iovdd out4_c out4 sg13g2_IOPadOut16mA
xp18 vss vdd vss iovdd out5_c out5 sg13g2_IOPadOut16mA
xp17 vss vdd vss iovdd out6_c out6 sg13g2_IOPadOut16mA
xp25 vss vdd vss iovdd sg13g2_IOPadVdd
xp16 vss vdd vss iovdd sg13g2_IOPadVss
xp27 vss vdd vss iovdd ck2_c ck2 sg13g2_IOPadIn
xp28 vss vdd vss iovdd ck3_c ck3 sg13g2_IOPadIn
xp29 vss vdd vss iovdd sg13g2_IOPadIOVdd
xp30 vss avdd vss avdd vldo net3 sg13g2_IOPadAnalog
xp31 vss avdd vss avdd vref vref_c sg13g2_IOPadAnalog
xp15 vss vdd vss iovdd ck6_c ck6 sg13g2_IOPadIn
xp14 vss vdd vss iovdd ck5_c ck5 sg13g2_IOPadIn
xp13 vss vdd vss iovdd ck4_c ck4 sg13g2_IOPadIn
xp12 vss vdd vss iovdd sg13g2_IOPadIOVss
xp11 vss vdd vss iovdd res_c res sg13g2_IOPadIn
xp10 vss avdd vss avdd sg13g2_IOPadVss
* noconn #net1
* noconn #net2
* noconn #net3
.ends

.GLOBAL GND
.GLOBAL VSS
.GLOBAL VDD
.end

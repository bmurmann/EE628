* Extracted by KLayout with SG13G2 LVS runset on : 03/05/2024 05:52

* cell sg13g2_RCClampInverter
* pin sub!
.SUBCKT sg13g2_RCClampInverter sub!
* device instance $1 r0 *1 7.72,6.54 sg13_hv_nmos
M$1 sub! \$3 sub! sub! sg13_hv_nmos W=125.99999999999999 L=9.499999999999996
* device instance $8 r0 *1 72.38,6.54 sg13_hv_nmos
M$8 sub! \$3 \$4 sub! sg13_hv_nmos W=107.99999999999999 L=0.4999999999999999
* device instance $27 r0 *1 18.44,29.91 sg13_hv_pmos
M$27 \$7 \$3 \$4 \$7 sg13_hv_pmos W=349.99999999999994 L=0.4999999999999999
.ENDS sg13g2_RCClampInverter

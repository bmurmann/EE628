.subckt RESISTOR in out
R1 in out 1k
.ends RESISTOR

.title KiCad schematic
.include "/home/maxwell/Desktop/ee699/sp-24-EE628/6_Test/2_PCB/test_board_1/TestBoardEDA/models/ADA4807-2.cir"

* voltage sources
V1 Net-_U1-VS+_ GND DC 5 
V2 GND Net-_U1-VS-_ DC 5 
V3 Net-_U1-IN1+_ GND DC 1 

XU1 Net-_U1-IN1+_ GND Net-_U1-VS+_ Net-_U1-VS-_ /out1 unconnected-_U1-IN2--Pad6_ ADA4807

.tran 1us 20ms
.print tran V(/out1)
.end


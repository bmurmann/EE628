** sch_path: /foss/designs/EE628/5_Design/3_Real_circuits/UHEE628_S2024.sch
.subckt UHEE628_S2024 vldo ck1 ck3 avdd ck2 VDD vref out1 in1 in2 out2 out3 in3 iovdd vhi vlo out4 in4 out5 in5 out6 in6 ck6 ck5
+ ck4 res VSS
*.PININFO in1:I in2:I in3:I in4:I in5:I in6:I iovdd:B vlo:B avdd:B out1:O out2:O out3:O out4:O out5:O out6:O VSS:B VDD:B vldo:B
*+ ck3:I ck2:I ck1:I vref:I res:I ck4:I ck5:I ck6:I vhi:B
x10 vref ck3 vldo ck1 ck2 ck1_c ck3_c net1 ck2_c out1_c in1 out1 in2 out2 out2_c in2_c VDD out3 in3_c in3 out3_c avdd iovdd vhi
+ vlo out4 in4_c in4 out4_c out5 in5_c out5_c in5 in6 in6_c out6 out6_c ck5_c ck4_c res_c ck6_c ck6 ck5 ck4 res in1_c VSS padring
x1 vhi vlo avdd VSS in1_c out1_c res_c ck1_c Team1
x2 vhi vlo avdd VSS in2_c out2_c res_c ck2_c template_idsm2
x4 vhi vlo avdd VSS in4_c out4_c res_c ck4_c template_idsm2
x5 vhi vlo avdd VSS in5_c out5_c res_c ck5_c Team5
* noconn #net1
x6 vhi vlo avdd VSS in6_c out6_c res_c ck6_c Team6
x7 vhi avdd res_c in3_c vlo out3_c VSS ck3_c Team3
.ends

* expanding   symbol:  padring.sym # of pins=47
** sym_path: /foss/designs/EE628/5_Design/3_Real_circuits/padring.sym
** sch_path: /foss/designs/EE628/5_Design/3_Real_circuits/padring.sch
.subckt padring vref ck3 vldo ck1 ck2 ck1_c ck3_c vref_c ck2_c out1_c in1 out1 in2 out2 out2_c in2_c vdd out3 in3_c in3 out3_c
+ avdd iovdd vhi vlo out4 in4_c in4 out4_c out5 in5_c out5_c in5 in6 in6_c out6 out6_c ck5_c ck4_c res_c ck6_c ck6 ck5 ck4 res in1_c vss
*.PININFO in1:I in2:I in3:I vhi:B vlo:B in4:I in5:I in6:I out1:O out2:O out3:O out4:O out5:O out6:O res:I ck4:I ck5:I ck6:I vref:I
*+ ck3:I ck2:I ck1:I in1_c:O in2_c:O in3_c:O in4_c:O in5_c:O in6_c:O res_c:O ck4_c:O ck5_c:O ck6_c:O out1_c:I out2_c:I out3_c:I out4_c:I
*+ out5_c:I out6_c:I vref_c:O ck3_c:O ck2_c:O ck1_c:O vldo:B avdd:B vss:B iovdd:B vdd:B
xp1 vss avdd vss avdd in1 in1_c sg13g2_IOPadAnalog
xp26 vss vdd vss iovdd ck1_c ck1 sg13g2_IOPadIn
xp24 vss vdd vss iovdd out1_c out1 sg13g2_IOPadOut16mA
xp32 vss avdd vss avdd sg13g2_IOPadVdd
xp9 vss avdd vss avdd sg13g2_IOPadVss
xp2 vss avdd vss avdd in2 in2_c sg13g2_IOPadAnalog
xp3 vss avdd vss avdd in3 in3_c sg13g2_IOPadAnalog
xp4 vss avdd vss avdd vhi net1 sg13g2_IOPadAnalog
xp5 vss avdd vss avdd vlo net2 sg13g2_IOPadAnalog
xp6 vss avdd vss avdd in4 in4_c sg13g2_IOPadAnalog
xp7 vss avdd vss avdd in5 in5_c sg13g2_IOPadAnalog
xp8 vss avdd vss avdd in6 in6_c sg13g2_IOPadAnalog
xp23 vss vdd vss iovdd out2_c out2 sg13g2_IOPadOut16mA
xp22 vss vdd vss iovdd out3_c out3 sg13g2_IOPadOut16mA
xp21 vss vdd vss iovdd sg13g2_IOPadIOVdd
xp20 vss vdd vss iovdd sg13g2_IOPadIOVss
xp19 vss vdd vss iovdd out4_c out4 sg13g2_IOPadOut16mA
xp18 vss vdd vss iovdd out5_c out5 sg13g2_IOPadOut16mA
xp17 vss vdd vss iovdd out6_c out6 sg13g2_IOPadOut16mA
xp25 vss vdd vss iovdd sg13g2_IOPadVdd
xp16 vss vdd vss iovdd sg13g2_IOPadVss
xp27 vss vdd vss iovdd ck2_c ck2 sg13g2_IOPadIn
xp28 vss vdd vss iovdd ck3_c ck3 sg13g2_IOPadIn
xp29 vss vdd vss iovdd sg13g2_IOPadIOVdd
xp30 vss avdd vss avdd vldo net3 sg13g2_IOPadAnalog
xp31 vss avdd vss avdd vref vref_c sg13g2_IOPadAnalog
xp15 vss vdd vss iovdd ck6_c ck6 sg13g2_IOPadIn
xp14 vss vdd vss iovdd ck5_c ck5 sg13g2_IOPadIn
xp13 vss vdd vss iovdd ck4_c ck4 sg13g2_IOPadIn
xp12 vss vdd vss iovdd sg13g2_IOPadIOVss
xp11 vss vdd vss iovdd res_c res sg13g2_IOPadIn
xp10 vss avdd vss avdd sg13g2_IOPadVss
* noconn #net1
* noconn #net2
* noconn #net3
.ends


* expanding   symbol:  /foss/designs/EE628/5_Design/3_Real_circuits/template_idsm2.sym # of pins=8
** sym_path: /foss/designs/EE628/5_Design/3_Real_circuits/template_idsm2.sym
** sch_path: /foss/designs/EE628/5_Design/3_Real_circuits/template_idsm2.sch
.subckt template_idsm2 vhi vlo vdda vssa vin dout res clkin
*.PININFO clkin:I res:I vin:I dout:O vssa:I vdda:I vlo:I vhi:I
x4 p1e p1 clkin p2 p2e template_clkgen
x1 res p1e p1 p2 vhi vdda vout1 vin vssa net1 vlo net3 template_stage
x2 res p2e p2 p1 vhi vdda vout2 vout1 vssa net2 vlo vmid2 template_stage
x3 vdda p2 net2 p1 net1 vout2 vmid2 vssa res dout template_comp
* noconn #net3
.ends


* expanding   symbol:  template_clkgen.sym # of pins=5
** sym_path: /foss/designs/EE628/5_Design/3_Real_circuits/template_clkgen.sym
** sch_path: /foss/designs/EE628/5_Design/3_Real_circuits/template_clkgen.sch
.subckt template_clkgen p1e p1 clkin p2 p2e
*.PININFO clkin:I p1e:O p1:O p2:O p2e:O
xn1 clkinbb b2 VDD VSS net11 sg13g2_nand2_2
xi7 net6 VDD VSS net9 sg13g2_inv_4
xi1 clkin VDD VSS clkinb sg13g2_inv_2
xi2 clkinb VDD VSS clkinbb sg13g2_inv_2
xn2 clkinb b1 VDD VSS net12 sg13g2_nand2_2
xi13 p1e VDD VSS b1 sg13g2_inv_4
xi8 net8 VDD VSS net10 sg13g2_inv_4
xi14 p2e VDD VSS b2 sg13g2_inv_4
xn3 a1 b1 VDD VSS net1 sg13g2_nand2_2
xn4 a2 b2 VDD VSS net3 sg13g2_nand2_2
xi11 a1 VDD VSS p1e sg13g2_inv_4
xi9 net9 VDD VSS a1 sg13g2_inv_4
x12 a2 VDD VSS p2e sg13g2_inv_4
xi10 net10 VDD VSS a2 sg13g2_inv_4
xi15 net1 VDD VSS net2 sg13g2_inv_4
xi17 net2 VDD VSS p1 sg13g2_inv_8
xi16 net3 VDD VSS net4 sg13g2_inv_4
xi18 net4 VDD VSS p2 sg13g2_inv_8
xi3 net11 VDD VSS net5 sg13g2_inv_4
xi5 net5 VDD VSS net6 sg13g2_inv_4
xi4 net12 VDD VSS net7 sg13g2_inv_4
xi6 net7 VDD VSS net8 sg13g2_inv_4
.ends


* expanding   symbol:  template_stage.sym # of pins=12
** sym_path: /foss/designs/EE628/5_Design/3_Real_circuits/template_stage.sym
** sch_path: /foss/designs/EE628/5_Design/3_Real_circuits/template_stage.sch
.subckt template_stage res pse ps pr vhi vdda vout vin vssa d vlo vmid
*.PININFO vout:O vdda:B res:I vin:I pse:I ps:I pr:I d:I vssa:B vhi:B vlo:B vmid:O
Mn vout vx3 vssa vssa sg13_lv_nmos L=1.5u W=2.5u ng=1 m=1
Mp vout vx3 vdda vdda sg13_lv_pmos L=1.5u W=10u ng=4 m=1
Mn3 vx1 gn vlo vssa sg13_lv_nmos L=0.13u W=0.5u ng=1 m=1
Mn4 vout res vx4 vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
x1 ps VDD VSS psb sg13g2_inv_1
Mp1 vx1 psb vin vdda sg13_lv_pmos L=0.13u W=6u ng=3 m=1
Mn5 vx1 ps vin vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
Mn1 vx4 pr vx2 vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
Mn2 vx4 ps vx3 vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
Mn6 vx2 pse vmid vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
Mn7 vmid vmid vssa vssa sg13_lv_nmos L=1.5u W=2.5u ng=1 m=1
Mp2 vmid vmid vdda vdda sg13_lv_pmos L=1.5u W=10u ng=4 m=1
x2 pr d VDD VSS gn sg13g2_and2_1
Mp3 vx1 gp vhi vdda sg13_lv_pmos L=0.13u W=1.5u ng=1 m=1
x3 d pr VDD VSS gp sg13g2_nand2b_1
C1 vx2 vx1 cap_cmim W=5.77e-6 L=5.77e-6 MF=1
C2 vx3 vx2 cap_cmim W=8.16e-6 L=8.16e-6 MF=1
C3 vx4 vout cap_cmim W=8.16e-6 L=8.16e-6 MF=1
.ends


* expanding   symbol:  template_comp.sym # of pins=10
** sym_path: /foss/designs/EE628/5_Design/3_Real_circuits/template_comp.sym
** sch_path: /foss/designs/EE628/5_Design/3_Real_circuits/template_comp.sch
.subckt template_comp vdda pc d ps dd vinm vinp vssa res dout
*.PININFO d:O pc:I vssa:B vdda:B ps:I res:I dd:O vinm:I vinp:I dout:O
M3m out1p out1m d2m vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M4m out1p out1m vdda vdda sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M5m out1p pc vdda vdda sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M2m d2m pc d1m vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M1m d1m vinm_samp vssa vssa sg13_lv_nmos L=1u W=2u ng=1 m=1
M3p out1m out1p d2p vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M4p out1m out1p vdda vdda sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M5p out1m pc vdda vdda sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M2p d2p pc d1p vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M1p d1p vinp vssa vssa sg13_lv_nmos L=1u W=2u ng=1 m=1
M32m dint net2 net1 VSS sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M2 dint net2 VDD VDD sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M3 dint out1m VDD VDD sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M21m net1 out1m VSS VSS sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M32p net2 dint net3 VSS sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M42p net2 dint VDD VDD sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M8 net2 out1p VDD VDD sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M21p net3 out1p VSS VSS sg13_lv_nmos L=0.13u W=2u ng=1 m=1
x1 ps dint dd net5 net4 VDD VSS sg13g2_dfrbp_2
x2 dint VDD VSS d sg13g2_buf_2
x3 res VDD VSS net4 sg13g2_inv_1
Mp1 vinm_samp psb vinm vdda sg13_lv_pmos L=0.13u W=6u ng=3 m=1
Mn5 vinm_samp ps vinm vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
C1 vinm_samp vssa cap_cmim W=5.77e-6 L=5.77e-6 MF=1
x4 ps VDD VSS psb sg13g2_inv_1
x5 dd VDD VSS dout sg13g2_inv_2
* noconn #net5
.ends

.GLOBAL VSS
.GLOBAL VDD
.end

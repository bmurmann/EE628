** sch_path: /foss/designs/EE628/5_Design/3_Real_circuits/UHEE628_S2024_top_schem.sch
.subckt UHEE628_S2024_top_schem in1 in2 in3 in4 in5 in6 iovdd vlo avdd out1 out2 out3 out4 out5 out6 VSS VDD vldo ck3 ck2 ck1 vref
+ res ck4 ck5 ck6 vhi
*.PININFO in1:I in2:I in3:I in4:I in5:I in6:I iovdd:B vlo:B avdd:B out1:O out2:O out3:O out4:O out5:O out6:O VSS:B VDD:B vldo:B
*+ ck3:I ck2:I ck1:I vref:I res:I ck4:I ck5:I ck6:I vhi:B
x10 vref ck3 vldo ck1 ck2 ck1_c ck3_c vref_c ck2_c out1_c in1 out1 in2 out2 out2_c in2_c VDD out3 in3_c in3 out3_c avdd iovdd vhi
+ vlo out4 in4_c in4 out4_c out5 in5_c out5_c in5 in6 in6_c out6 out6_c ck5_c ck4_c res_c ck6_c ck6 ck5 ck4 res in1_c VSS padring
x1 vhi vlo avdd VSS in1_c out1_c res_c ck1_c IDSM2_t1
x2 vlo vhi vldo VSS iovdd vref_c in2_c out2_c res_c ck2_c Team_2
x4 vhi vlo avdd VSS in4_c out4_c res_c ck4_c IDSM2_T4
x5 vhi vlo out5_c avdd VSS in5_c res_c ck5_c Team5
x6 vhi vlo avdd VSS in6_c out6_c res_c ck6_c Team6_inner
x3 vhi vlo avdd VSS in3_c out3_c res_c ck3_c Team3
.ends

* expanding   symbol:  padring.sym # of pins=47
** sym_path: /foss/designs/EE628/5_Design/3_Real_circuits/padring.sym
** sch_path: /foss/designs/EE628/5_Design/3_Real_circuits/padring.sch
.subckt padring vref ck3 vldo ck1 ck2 ck1_c ck3_c vref_c ck2_c out1_c in1 out1 in2 out2 out2_c in2_c vdd out3 in3_c in3 out3_c
+ avdd iovdd vhi vlo out4 in4_c in4 out4_c out5 in5_c out5_c in5 in6 in6_c out6 out6_c ck5_c ck4_c res_c ck6_c ck6 ck5 ck4 res in1_c vss
*.PININFO in1:I in2:I in3:I vhi:B vlo:B in4:I in5:I in6:I out1:O out2:O out3:O out4:O out5:O out6:O res:I ck4:I ck5:I ck6:I vref:I
*+ ck3:I ck2:I ck1:I in1_c:O in2_c:O in3_c:O in4_c:O in5_c:O in6_c:O res_c:O ck4_c:O ck5_c:O ck6_c:O out1_c:I out2_c:I out3_c:I out4_c:I
*+ out5_c:I out6_c:I vref_c:O ck3_c:O ck2_c:O ck1_c:O vldo:B avdd:B vss:B iovdd:B vdd:B
xp1 vss avdd vss avdd in1 in1_c sg13g2_IOPadAnalog
xp26 vss vdd vss iovdd ck1_c ck1 sg13g2_IOPadIn
xp24 vss vdd vss iovdd out1_c out1 sg13g2_IOPadOut16mA
xp32 vss avdd vss avdd sg13g2_IOPadVdd
xp9 vss avdd vss avdd sg13g2_IOPadVss
xp2 vss avdd vss avdd in2 in2_c sg13g2_IOPadAnalog
xp3 vss avdd vss avdd in3 in3_c sg13g2_IOPadAnalog
xp4 vss avdd vss avdd vhi net1 sg13g2_IOPadAnalog
xp5 vss avdd vss avdd vlo net2 sg13g2_IOPadAnalog
xp6 vss avdd vss avdd in4 in4_c sg13g2_IOPadAnalog
xp7 vss avdd vss avdd in5 in5_c sg13g2_IOPadAnalog
xp8 vss avdd vss avdd in6 in6_c sg13g2_IOPadAnalog
xp23 vss vdd vss iovdd out2_c out2 sg13g2_IOPadOut16mA
xp22 vss vdd vss iovdd out3_c out3 sg13g2_IOPadOut16mA
xp21 vss vdd vss iovdd sg13g2_IOPadIOVdd
xp20 vss vdd vss iovdd sg13g2_IOPadIOVss
xp19 vss vdd vss iovdd out4_c out4 sg13g2_IOPadOut16mA
xp18 vss vdd vss iovdd out5_c out5 sg13g2_IOPadOut16mA
xp17 vss vdd vss iovdd out6_c out6 sg13g2_IOPadOut16mA
xp25 vss vdd vss iovdd sg13g2_IOPadVdd
xp16 vss vdd vss iovdd sg13g2_IOPadVss
xp27 vss vdd vss iovdd ck2_c ck2 sg13g2_IOPadIn
xp28 vss vdd vss iovdd ck3_c ck3 sg13g2_IOPadIn
xp29 vss vdd vss iovdd sg13g2_IOPadIOVdd
xp30 vss avdd vss avdd vldo net3 sg13g2_IOPadAnalog
xp31 vss avdd vss avdd vref vref_c sg13g2_IOPadAnalog
xp15 vss vdd vss iovdd ck6_c ck6 sg13g2_IOPadIn
xp14 vss vdd vss iovdd ck5_c ck5 sg13g2_IOPadIn
xp13 vss vdd vss iovdd ck4_c ck4 sg13g2_IOPadIn
xp12 vss vdd vss iovdd sg13g2_IOPadIOVss
xp11 vss vdd vss iovdd res_c res sg13g2_IOPadIn
xp10 vss avdd vss avdd sg13g2_IOPadVss
* noconn #net1
* noconn #net2
* noconn #net3
.ends


* expanding   symbol:  /foss/designs/EE628/5_Design/4_Layout/Team 5/Team5.sym # of pins=8
** sym_path: /foss/designs/EE628/5_Design/4_Layout/Team 5/Team5.sym
** sch_path: /foss/designs/EE628/5_Design/4_Layout/Team 5/Team5.sch
.subckt Team5 vhi vlo dd vdda vssa vin res clkin
*.PININFO vhi:I vlo:I vdda:I vssa:I vin:I res:I dd:O clkin:I
*  x2 -  Team5_split1  IS MISSING !!!!
*  x1 -  Team5_split2  IS MISSING !!!!
.ends

.GLOBAL VSS
.GLOBAL VDD
.end

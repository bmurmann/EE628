* Extracted by KLayout with SG13G2 LVS runset on : 09/05/2024 23:30

* cell clock_5_splitTop
* pin inv_bottom
* pin VDD
* pin clkin
* pin nand_B2
* pin VSS
.SUBCKT clock_5_splitTop inv_bottom VDD clkin nand_B2 VSS
* device instance $1 r0 *1 5.9,-6.712 sg13_lv_nmos
M$1 \$3 nand_B2 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $3 r0 *1 6.93,-6.712 sg13_lv_nmos
M$3 \$3 \$69 \$15 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $5 r0 *1 31.086,-6.712 sg13_lv_nmos
M$5 \$4 \$21 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $7 r0 *1 32.116,-6.712 sg13_lv_nmos
M$7 \$4 \$19 \$22 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $9 r0 *1 9.164,-6.687 sg13_lv_nmos
M$9 VSS \$15 \$16 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $13 r0 *1 12.579,-6.687 sg13_lv_nmos
M$13 VSS \$16 \$17 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $17 r0 *1 15.815,-6.687 sg13_lv_nmos
M$17 VSS \$17 \$18 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $21 r0 *1 19.34,-6.687 sg13_lv_nmos
M$21 VSS \$18 \$19 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $25 r0 *1 23.197,-6.687 sg13_lv_nmos
M$25 VSS \$19 inv_bottom VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $29 r0 *1 27.166,-6.687 sg13_lv_nmos
M$29 VSS inv_bottom \$21 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $33 r0 *1 34.77,-6.687 sg13_lv_nmos
M$33 VSS \$22 \$23 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $37 r0 *1 38.166,-6.687 sg13_lv_nmos
M$37 VSS \$23 \$24 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $45 r0 *1 0.011,1.281 sg13_lv_nmos
M$45 VSS clkin nand_B2 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $47 r0 *1 2.532,1.281 sg13_lv_nmos
M$47 VSS nand_B2 \$86 VSS sg13_lv_nmos W=1.48 L=0.13
* device instance $49 r0 *1 5.178,1.256 sg13_lv_nmos
M$49 \$63 \$86 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $51 r0 *1 6.208,1.256 sg13_lv_nmos
M$51 \$63 \$21 \$87 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $53 r0 *1 8.541,1.282 sg13_lv_nmos
M$53 VSS \$87 \$64 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $57 r0 *1 13.009,1.282 sg13_lv_nmos
M$57 VSS \$64 \$65 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $61 r0 *1 16.425,1.282 sg13_lv_nmos
M$61 VSS \$65 \$66 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $65 r0 *1 19.945,1.282 sg13_lv_nmos
M$65 VSS \$66 \$67 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $69 r0 *1 23.802,1.282 sg13_lv_nmos
M$69 VSS \$67 \$68 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $73 r0 *1 27.771,1.282 sg13_lv_nmos
M$73 VSS \$68 \$69 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $77 r0 *1 31.441,1.257 sg13_lv_nmos
M$77 \$70 \$69 VSS VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $79 r0 *1 32.471,1.257 sg13_lv_nmos
M$79 \$70 \$67 \$88 VSS sg13_lv_nmos W=1.44 L=0.13
* device instance $81 r0 *1 35.125,1.282 sg13_lv_nmos
M$81 VSS \$88 \$71 VSS sg13_lv_nmos W=2.96 L=0.13
* device instance $85 r0 *1 38.521,1.282 sg13_lv_nmos
M$85 VSS \$71 \$89 VSS sg13_lv_nmos W=5.920000000000001 L=0.13
* device instance $93 r0 *1 5.9,-5.027 sg13_lv_pmos
M$93 VDD nand_B2 \$15 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $95 r0 *1 6.93,-5.027 sg13_lv_pmos
M$95 VDD \$69 \$15 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $97 r0 *1 9.164,-5.027 sg13_lv_pmos
M$97 VDD \$15 \$16 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $101 r0 *1 12.579,-5.027 sg13_lv_pmos
M$101 VDD \$16 \$17 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $105 r0 *1 15.815,-5.027 sg13_lv_pmos
M$105 VDD \$17 \$18 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $109 r0 *1 19.34,-5.027 sg13_lv_pmos
M$109 VDD \$18 \$19 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $113 r0 *1 23.197,-5.027 sg13_lv_pmos
M$113 VDD \$19 inv_bottom VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $117 r0 *1 27.166,-5.027 sg13_lv_pmos
M$117 VDD inv_bottom \$21 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $121 r0 *1 31.086,-5.027 sg13_lv_pmos
M$121 VDD \$21 \$22 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $123 r0 *1 32.116,-5.027 sg13_lv_pmos
M$123 VDD \$19 \$22 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $125 r0 *1 34.77,-5.027 sg13_lv_pmos
M$125 VDD \$22 \$23 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $129 r0 *1 38.166,-5.027 sg13_lv_pmos
M$129 VDD \$23 \$24 VDD sg13_lv_pmos W=8.96 L=0.13
* device instance $137 r0 *1 0.001,2.941 sg13_lv_pmos
M$137 VDD clkin nand_B2 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $139 r0 *1 2.522,2.941 sg13_lv_pmos
M$139 VDD nand_B2 \$86 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $141 r0 *1 5.178,2.941 sg13_lv_pmos
M$141 VDD \$86 \$87 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $143 r0 *1 6.208,2.941 sg13_lv_pmos
M$143 VDD \$21 \$87 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $145 r0 *1 8.541,2.942 sg13_lv_pmos
M$145 VDD \$87 \$64 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $149 r0 *1 13.009,2.942 sg13_lv_pmos
M$149 VDD \$64 \$65 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $153 r0 *1 16.425,2.942 sg13_lv_pmos
M$153 VDD \$65 \$66 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $157 r0 *1 19.945,2.942 sg13_lv_pmos
M$157 VDD \$66 \$67 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $161 r0 *1 23.802,2.942 sg13_lv_pmos
M$161 VDD \$67 \$68 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $165 r0 *1 27.771,2.942 sg13_lv_pmos
M$165 VDD \$68 \$69 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $169 r0 *1 31.441,2.942 sg13_lv_pmos
M$169 VDD \$69 \$88 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $171 r0 *1 32.471,2.942 sg13_lv_pmos
M$171 VDD \$67 \$88 VDD sg13_lv_pmos W=2.24 L=0.13
* device instance $173 r0 *1 35.125,2.942 sg13_lv_pmos
M$173 VDD \$88 \$71 VDD sg13_lv_pmos W=4.48 L=0.13
* device instance $177 r0 *1 38.521,2.942 sg13_lv_pmos
M$177 VDD \$71 \$89 VDD sg13_lv_pmos W=8.96 L=0.13
.ENDS clock_5_splitTop
